

logic [15:0] PLUT [32] = '{
    16'h10c5,
    16'h0,
    16'h10c4,
    16'h882,
    16'hca4,
    16'h460,
    16'h420,
    16'h20,
    16'h862,
    16'h421,
    16'h861,
    16'h441,
    16'h41,
    16'h8a2,
    16'h881,
    16'h440,
    16'h8a1,
    16'h8c1,
    16'hcc1,
    16'hcc2,
    16'h480,
    16'hcc3,
    16'h8a0,
    16'h10c3,
    16'h14e5,
    16'h10e4,
    16'hffff,
    16'hffff,
    16'hffff,
    16'hffff,
    16'hffff,
    16'hffff
};

task automatic setup_cel_core(ref McoreRegs_t mcoreClass);
/*Cel Vars setup begin*/
    mcoreClass.set_cel_int_var(HDDX1616_ID, 32'h0);
    mcoreClass.set_cel_int_var(HDDY1616_ID, 32'h0);
    mcoreClass.set_cel_int_var(HDX1616_ID, 32'h10000);
    mcoreClass.set_cel_int_var(HDY1616_ID, 32'h0);
    mcoreClass.set_cel_int_var(VDX1616_ID, 32'h0);
    mcoreClass.set_cel_int_var(VDY1616_ID, 32'h10000);
    mcoreClass.set_cel_int_var(XPOS1616_ID, 32'h1349000);
    mcoreClass.set_cel_int_var(YPOS1616_ID, 32'h6a0000);
    mcoreClass.set_cel_int_var(HDX1616_2_ID, 32'h0);
    mcoreClass.set_cel_int_var(HDY1616_2_ID, 32'h0);
    mcoreClass.set_cel_int_var(TEXTURE_WI_START_ID, 32'h0);
    mcoreClass.set_cel_int_var(TEXTURE_HI_START_ID, 32'h0);
    mcoreClass.set_cel_int_var(TEXEL_INCX_ID, 32'h1);
    mcoreClass.set_cel_int_var(TEXEL_INCY_ID, 32'h1);
    mcoreClass.set_cel_int_var(TEXTURE_WI_LIM_ID, 32'h56);
    mcoreClass.set_cel_int_var(TEXTURE_HI_LIM_ID, 32'hb0);
    mcoreClass.set_cel_int_var(TEXEL_FUN_NUMBER_ID, 32'h1);
    mcoreClass.set_cel_int_var(SPRWI_ID, 32'h2);
    mcoreClass.set_cel_int_var(SPRHI_ID, 32'h16);
    mcoreClass.set_cel_int_var(BITCALC_ID, 32'h180);
    mcoreClass.set_cel_uint_var(BITADDR_ID, 32'h0);
    mcoreClass.set_cel_uint_var(BITBUFLEN_ID, 32'h0);
    mcoreClass.set_cel_uint_var(BITBUF_ID, 32'h0);
    mcoreClass.set_cel_uint_var(CCBFLAGS_ID, 32'h3fbec000);
    mcoreClass.set_cel_uint_var(PIXC_ID, 32'h1f811f00);
    mcoreClass.set_cel_uint_var(PRE0_ID, 32'h544);
    mcoreClass.set_cel_uint_var(PRE1_ID, 32'h1001);
    mcoreClass.set_cel_uint_var(TARGETPROJ_ID, 32'h0);
    mcoreClass.set_cel_uint_var(SRCDATA_ID, 32'h0);
    mcoreClass.set_cel_uint_var(PLUTF_ID, 32'h0);
    mcoreClass.set_cel_uint_var(PDATF_ID, 32'h0);
    mcoreClass.set_cel_uint_var(NCCBF_ID, 32'h0);
    mcoreClass.set_cel_uint_var(PXOR1_ID, 32'hffffffff);
    mcoreClass.set_cel_uint_var(PXOR2_ID, 32'h0);
/*Cel Vars setup end*/


/*Setup mregs begin*/
    mcoreClass.set_mregs(32'h0, 32'h1020000);
    mcoreClass.set_mregs(32'h1, 32'h0);
    mcoreClass.set_mregs(32'h2, 32'h0);
    mcoreClass.set_mregs(32'h3, 32'h0);
    mcoreClass.set_mregs(32'h4, 32'h29);
    mcoreClass.set_mregs(32'h5, 32'h0);
    mcoreClass.set_mregs(32'h6, 32'h0);
    mcoreClass.set_mregs(32'h7, 32'h0);
    mcoreClass.set_mregs(32'h8, 32'hffef7fff);
    mcoreClass.set_mregs(32'h9, 32'h0);
    mcoreClass.set_mregs(32'ha, 32'h0);
    mcoreClass.set_mregs(32'hb, 32'h0);
    mcoreClass.set_mregs(32'hc, 32'h0);
    mcoreClass.set_mregs(32'hd, 32'h0);
    mcoreClass.set_mregs(32'he, 32'h0);
    mcoreClass.set_mregs(32'hf, 32'h0);
    mcoreClass.set_mregs(32'h10, 32'h0);
    mcoreClass.set_mregs(32'h11, 32'h0);
    mcoreClass.set_mregs(32'h12, 32'h0);
    mcoreClass.set_mregs(32'h13, 32'h0);
    mcoreClass.set_mregs(32'h14, 32'h0);
    mcoreClass.set_mregs(32'h15, 32'h0);
    mcoreClass.set_mregs(32'h16, 32'h0);
    mcoreClass.set_mregs(32'h17, 32'h0);
    mcoreClass.set_mregs(32'h18, 32'h0);
    mcoreClass.set_mregs(32'h19, 32'h0);
    mcoreClass.set_mregs(32'h1a, 32'h0);
    mcoreClass.set_mregs(32'h1b, 32'h0);
    mcoreClass.set_mregs(32'h1c, 32'h0);
    mcoreClass.set_mregs(32'h1d, 32'h0);
    mcoreClass.set_mregs(32'h1e, 32'h0);
    mcoreClass.set_mregs(32'h1f, 32'h0);
    mcoreClass.set_mregs(32'h20, 32'h0);
    mcoreClass.set_mregs(32'h21, 32'h0);
    mcoreClass.set_mregs(32'h22, 32'h0);
    mcoreClass.set_mregs(32'h23, 32'h0);
    mcoreClass.set_mregs(32'h24, 32'h0);
    mcoreClass.set_mregs(32'h25, 32'h0);
    mcoreClass.set_mregs(32'h26, 32'h0);
    mcoreClass.set_mregs(32'h27, 32'h0);
    mcoreClass.set_mregs(32'h28, 32'h10);
    mcoreClass.set_mregs(32'h29, 32'h0);
    mcoreClass.set_mregs(32'h2a, 32'h0);
    mcoreClass.set_mregs(32'h2b, 32'h0);
    mcoreClass.set_mregs(32'h2c, 32'h0);
    mcoreClass.set_mregs(32'h2d, 32'h0);
    mcoreClass.set_mregs(32'h2e, 32'h0);
    mcoreClass.set_mregs(32'h2f, 32'h0);
    mcoreClass.set_mregs(32'h30, 32'h0);
    mcoreClass.set_mregs(32'h31, 32'h0);
    mcoreClass.set_mregs(32'h32, 32'h0);
    mcoreClass.set_mregs(32'h33, 32'h0);
    mcoreClass.set_mregs(32'h34, 32'h0);
    mcoreClass.set_mregs(32'h35, 32'h0);
    mcoreClass.set_mregs(32'h36, 32'h0);
    mcoreClass.set_mregs(32'h37, 32'h0);
    mcoreClass.set_mregs(32'h38, 32'h0);
    mcoreClass.set_mregs(32'h39, 32'h0);
    mcoreClass.set_mregs(32'h3a, 32'h0);
    mcoreClass.set_mregs(32'h3b, 32'h0);
    mcoreClass.set_mregs(32'h3c, 32'h0);
    mcoreClass.set_mregs(32'h3d, 32'h0);
    mcoreClass.set_mregs(32'h3e, 32'h0);
    mcoreClass.set_mregs(32'h3f, 32'h0);
    mcoreClass.set_mregs(32'h40, 32'h0);
    mcoreClass.set_mregs(32'h41, 32'h0);
    mcoreClass.set_mregs(32'h42, 32'h0);
    mcoreClass.set_mregs(32'h43, 32'h0);
    mcoreClass.set_mregs(32'h44, 32'h0);
    mcoreClass.set_mregs(32'h45, 32'h0);
    mcoreClass.set_mregs(32'h46, 32'h0);
    mcoreClass.set_mregs(32'h47, 32'h0);
    mcoreClass.set_mregs(32'h48, 32'h0);
    mcoreClass.set_mregs(32'h49, 32'h0);
    mcoreClass.set_mregs(32'h4a, 32'h0);
    mcoreClass.set_mregs(32'h4b, 32'h0);
    mcoreClass.set_mregs(32'h4c, 32'h0);
    mcoreClass.set_mregs(32'h4d, 32'h0);
    mcoreClass.set_mregs(32'h4e, 32'h0);
    mcoreClass.set_mregs(32'h4f, 32'h0);
    mcoreClass.set_mregs(32'h50, 32'h0);
    mcoreClass.set_mregs(32'h51, 32'h0);
    mcoreClass.set_mregs(32'h52, 32'h0);
    mcoreClass.set_mregs(32'h53, 32'h0);
    mcoreClass.set_mregs(32'h54, 32'h0);
    mcoreClass.set_mregs(32'h55, 32'h0);
    mcoreClass.set_mregs(32'h56, 32'h0);
    mcoreClass.set_mregs(32'h57, 32'h0);
    mcoreClass.set_mregs(32'h58, 32'h0);
    mcoreClass.set_mregs(32'h59, 32'h0);
    mcoreClass.set_mregs(32'h5a, 32'h0);
    mcoreClass.set_mregs(32'h5b, 32'h0);
    mcoreClass.set_mregs(32'h5c, 32'h0);
    mcoreClass.set_mregs(32'h5d, 32'h0);
    mcoreClass.set_mregs(32'h5e, 32'h0);
    mcoreClass.set_mregs(32'h5f, 32'h0);
    mcoreClass.set_mregs(32'h60, 32'h0);
    mcoreClass.set_mregs(32'h61, 32'h0);
    mcoreClass.set_mregs(32'h62, 32'h0);
    mcoreClass.set_mregs(32'h63, 32'h0);
    mcoreClass.set_mregs(32'h64, 32'h0);
    mcoreClass.set_mregs(32'h65, 32'h0);
    mcoreClass.set_mregs(32'h66, 32'h0);
    mcoreClass.set_mregs(32'h67, 32'h0);
    mcoreClass.set_mregs(32'h68, 32'h0);
    mcoreClass.set_mregs(32'h69, 32'h0);
    mcoreClass.set_mregs(32'h6a, 32'h0);
    mcoreClass.set_mregs(32'h6b, 32'h0);
    mcoreClass.set_mregs(32'h6c, 32'h0);
    mcoreClass.set_mregs(32'h6d, 32'h0);
    mcoreClass.set_mregs(32'h6e, 32'h0);
    mcoreClass.set_mregs(32'h6f, 32'h0);
    mcoreClass.set_mregs(32'h70, 32'h0);
    mcoreClass.set_mregs(32'h71, 32'h0);
    mcoreClass.set_mregs(32'h72, 32'h0);
    mcoreClass.set_mregs(32'h73, 32'h0);
    mcoreClass.set_mregs(32'h74, 32'h0);
    mcoreClass.set_mregs(32'h75, 32'h0);
    mcoreClass.set_mregs(32'h76, 32'h0);
    mcoreClass.set_mregs(32'h77, 32'h0);
    mcoreClass.set_mregs(32'h78, 32'h0);
    mcoreClass.set_mregs(32'h79, 32'h0);
    mcoreClass.set_mregs(32'h7a, 32'h0);
    mcoreClass.set_mregs(32'h7b, 32'h0);
    mcoreClass.set_mregs(32'h7c, 32'h0);
    mcoreClass.set_mregs(32'h7d, 32'h0);
    mcoreClass.set_mregs(32'h7e, 32'h0);
    mcoreClass.set_mregs(32'h7f, 32'h0);
    mcoreClass.set_mregs(32'h80, 32'h0);
    mcoreClass.set_mregs(32'h81, 32'h0);
    mcoreClass.set_mregs(32'h82, 32'h0);
    mcoreClass.set_mregs(32'h83, 32'h0);
    mcoreClass.set_mregs(32'h84, 32'h0);
    mcoreClass.set_mregs(32'h85, 32'h0);
    mcoreClass.set_mregs(32'h86, 32'h0);
    mcoreClass.set_mregs(32'h87, 32'h0);
    mcoreClass.set_mregs(32'h88, 32'h0);
    mcoreClass.set_mregs(32'h89, 32'h0);
    mcoreClass.set_mregs(32'h8a, 32'h0);
    mcoreClass.set_mregs(32'h8b, 32'h0);
    mcoreClass.set_mregs(32'h8c, 32'h0);
    mcoreClass.set_mregs(32'h8d, 32'h0);
    mcoreClass.set_mregs(32'h8e, 32'h0);
    mcoreClass.set_mregs(32'h8f, 32'h0);
    mcoreClass.set_mregs(32'h90, 32'h0);
    mcoreClass.set_mregs(32'h91, 32'h0);
    mcoreClass.set_mregs(32'h92, 32'h0);
    mcoreClass.set_mregs(32'h93, 32'h0);
    mcoreClass.set_mregs(32'h94, 32'h0);
    mcoreClass.set_mregs(32'h95, 32'h0);
    mcoreClass.set_mregs(32'h96, 32'h0);
    mcoreClass.set_mregs(32'h97, 32'h0);
    mcoreClass.set_mregs(32'h98, 32'h0);
    mcoreClass.set_mregs(32'h99, 32'h0);
    mcoreClass.set_mregs(32'h9a, 32'h0);
    mcoreClass.set_mregs(32'h9b, 32'h0);
    mcoreClass.set_mregs(32'h9c, 32'h0);
    mcoreClass.set_mregs(32'h9d, 32'h0);
    mcoreClass.set_mregs(32'h9e, 32'h0);
    mcoreClass.set_mregs(32'h9f, 32'h0);
    mcoreClass.set_mregs(32'ha0, 32'h0);
    mcoreClass.set_mregs(32'ha1, 32'h0);
    mcoreClass.set_mregs(32'ha2, 32'h0);
    mcoreClass.set_mregs(32'ha3, 32'h0);
    mcoreClass.set_mregs(32'ha4, 32'h0);
    mcoreClass.set_mregs(32'ha5, 32'h0);
    mcoreClass.set_mregs(32'ha6, 32'h0);
    mcoreClass.set_mregs(32'ha7, 32'h0);
    mcoreClass.set_mregs(32'ha8, 32'h0);
    mcoreClass.set_mregs(32'ha9, 32'h0);
    mcoreClass.set_mregs(32'haa, 32'h0);
    mcoreClass.set_mregs(32'hab, 32'h0);
    mcoreClass.set_mregs(32'hac, 32'h0);
    mcoreClass.set_mregs(32'had, 32'h0);
    mcoreClass.set_mregs(32'hae, 32'h0);
    mcoreClass.set_mregs(32'haf, 32'h0);
    mcoreClass.set_mregs(32'hb0, 32'h0);
    mcoreClass.set_mregs(32'hb1, 32'h0);
    mcoreClass.set_mregs(32'hb2, 32'h0);
    mcoreClass.set_mregs(32'hb3, 32'h0);
    mcoreClass.set_mregs(32'hb4, 32'h0);
    mcoreClass.set_mregs(32'hb5, 32'h0);
    mcoreClass.set_mregs(32'hb6, 32'h0);
    mcoreClass.set_mregs(32'hb7, 32'h0);
    mcoreClass.set_mregs(32'hb8, 32'h0);
    mcoreClass.set_mregs(32'hb9, 32'h0);
    mcoreClass.set_mregs(32'hba, 32'h0);
    mcoreClass.set_mregs(32'hbb, 32'h0);
    mcoreClass.set_mregs(32'hbc, 32'h0);
    mcoreClass.set_mregs(32'hbd, 32'h0);
    mcoreClass.set_mregs(32'hbe, 32'h0);
    mcoreClass.set_mregs(32'hbf, 32'h0);
    mcoreClass.set_mregs(32'hc0, 32'h0);
    mcoreClass.set_mregs(32'hc1, 32'h0);
    mcoreClass.set_mregs(32'hc2, 32'h0);
    mcoreClass.set_mregs(32'hc3, 32'h0);
    mcoreClass.set_mregs(32'hc4, 32'h0);
    mcoreClass.set_mregs(32'hc5, 32'h0);
    mcoreClass.set_mregs(32'hc6, 32'h0);
    mcoreClass.set_mregs(32'hc7, 32'h0);
    mcoreClass.set_mregs(32'hc8, 32'h0);
    mcoreClass.set_mregs(32'hc9, 32'h0);
    mcoreClass.set_mregs(32'hca, 32'h0);
    mcoreClass.set_mregs(32'hcb, 32'h0);
    mcoreClass.set_mregs(32'hcc, 32'h0);
    mcoreClass.set_mregs(32'hcd, 32'h0);
    mcoreClass.set_mregs(32'hce, 32'h0);
    mcoreClass.set_mregs(32'hcf, 32'h0);
    mcoreClass.set_mregs(32'hd0, 32'h0);
    mcoreClass.set_mregs(32'hd1, 32'h0);
    mcoreClass.set_mregs(32'hd2, 32'h0);
    mcoreClass.set_mregs(32'hd3, 32'h0);
    mcoreClass.set_mregs(32'hd4, 32'h0);
    mcoreClass.set_mregs(32'hd5, 32'h0);
    mcoreClass.set_mregs(32'hd6, 32'h0);
    mcoreClass.set_mregs(32'hd7, 32'h0);
    mcoreClass.set_mregs(32'hd8, 32'h0);
    mcoreClass.set_mregs(32'hd9, 32'h0);
    mcoreClass.set_mregs(32'hda, 32'h0);
    mcoreClass.set_mregs(32'hdb, 32'h0);
    mcoreClass.set_mregs(32'hdc, 32'h0);
    mcoreClass.set_mregs(32'hdd, 32'h0);
    mcoreClass.set_mregs(32'hde, 32'h0);
    mcoreClass.set_mregs(32'hdf, 32'h0);
    mcoreClass.set_mregs(32'he0, 32'h0);
    mcoreClass.set_mregs(32'he1, 32'h0);
    mcoreClass.set_mregs(32'he2, 32'h0);
    mcoreClass.set_mregs(32'he3, 32'h0);
    mcoreClass.set_mregs(32'he4, 32'h0);
    mcoreClass.set_mregs(32'he5, 32'h0);
    mcoreClass.set_mregs(32'he6, 32'h0);
    mcoreClass.set_mregs(32'he7, 32'h0);
    mcoreClass.set_mregs(32'he8, 32'h0);
    mcoreClass.set_mregs(32'he9, 32'h0);
    mcoreClass.set_mregs(32'hea, 32'h0);
    mcoreClass.set_mregs(32'heb, 32'h0);
    mcoreClass.set_mregs(32'hec, 32'h0);
    mcoreClass.set_mregs(32'hed, 32'h0);
    mcoreClass.set_mregs(32'hee, 32'h0);
    mcoreClass.set_mregs(32'hef, 32'h0);
    mcoreClass.set_mregs(32'hf0, 32'h0);
    mcoreClass.set_mregs(32'hf1, 32'h0);
    mcoreClass.set_mregs(32'hf2, 32'h0);
    mcoreClass.set_mregs(32'hf3, 32'h0);
    mcoreClass.set_mregs(32'hf4, 32'h0);
    mcoreClass.set_mregs(32'hf5, 32'h0);
    mcoreClass.set_mregs(32'hf6, 32'h0);
    mcoreClass.set_mregs(32'hf7, 32'h0);
    mcoreClass.set_mregs(32'hf8, 32'h0);
    mcoreClass.set_mregs(32'hf9, 32'h0);
    mcoreClass.set_mregs(32'hfa, 32'h0);
    mcoreClass.set_mregs(32'hfb, 32'h0);
    mcoreClass.set_mregs(32'hfc, 32'h0);
    mcoreClass.set_mregs(32'hfd, 32'h0);
    mcoreClass.set_mregs(32'hfe, 32'h0);
    mcoreClass.set_mregs(32'hff, 32'h0);
    mcoreClass.set_mregs(32'h100, 32'h0);
    mcoreClass.set_mregs(32'h101, 32'h0);
    mcoreClass.set_mregs(32'h102, 32'h0);
    mcoreClass.set_mregs(32'h103, 32'h0);
    mcoreClass.set_mregs(32'h104, 32'h0);
    mcoreClass.set_mregs(32'h105, 32'h0);
    mcoreClass.set_mregs(32'h106, 32'h0);
    mcoreClass.set_mregs(32'h107, 32'h0);
    mcoreClass.set_mregs(32'h108, 32'h0);
    mcoreClass.set_mregs(32'h109, 32'h0);
    mcoreClass.set_mregs(32'h10a, 32'h0);
    mcoreClass.set_mregs(32'h10b, 32'h0);
    mcoreClass.set_mregs(32'h10c, 32'h0);
    mcoreClass.set_mregs(32'h10d, 32'h0);
    mcoreClass.set_mregs(32'h10e, 32'h0);
    mcoreClass.set_mregs(32'h10f, 32'h0);
    mcoreClass.set_mregs(32'h110, 32'he1500000);
    mcoreClass.set_mregs(32'h111, 32'h0);
    mcoreClass.set_mregs(32'h112, 32'h0);
    mcoreClass.set_mregs(32'h113, 32'h0);
    mcoreClass.set_mregs(32'h114, 32'h0);
    mcoreClass.set_mregs(32'h115, 32'h0);
    mcoreClass.set_mregs(32'h116, 32'h0);
    mcoreClass.set_mregs(32'h117, 32'h0);
    mcoreClass.set_mregs(32'h118, 32'h0);
    mcoreClass.set_mregs(32'h119, 32'h0);
    mcoreClass.set_mregs(32'h11a, 32'h0);
    mcoreClass.set_mregs(32'h11b, 32'h0);
    mcoreClass.set_mregs(32'h11c, 32'h0);
    mcoreClass.set_mregs(32'h11d, 32'h0);
    mcoreClass.set_mregs(32'h11e, 32'h0);
    mcoreClass.set_mregs(32'h11f, 32'h0);
    mcoreClass.set_mregs(32'h120, 32'h0);
    mcoreClass.set_mregs(32'h121, 32'h0);
    mcoreClass.set_mregs(32'h122, 32'h0);
    mcoreClass.set_mregs(32'h123, 32'h0);
    mcoreClass.set_mregs(32'h124, 32'h0);
    mcoreClass.set_mregs(32'h125, 32'h0);
    mcoreClass.set_mregs(32'h126, 32'h0);
    mcoreClass.set_mregs(32'h127, 32'h0);
    mcoreClass.set_mregs(32'h128, 32'h0);
    mcoreClass.set_mregs(32'h129, 32'h0);
    mcoreClass.set_mregs(32'h12a, 32'h0);
    mcoreClass.set_mregs(32'h12b, 32'h0);
    mcoreClass.set_mregs(32'h12c, 32'h0);
    mcoreClass.set_mregs(32'h12d, 32'h0);
    mcoreClass.set_mregs(32'h12e, 32'h0);
    mcoreClass.set_mregs(32'h12f, 32'h0);
    mcoreClass.set_mregs(32'h130, 32'h1414);
    mcoreClass.set_mregs(32'h131, 32'h0);
    mcoreClass.set_mregs(32'h132, 32'h0);
    mcoreClass.set_mregs(32'h133, 32'h0);
    mcoreClass.set_mregs(32'h134, 32'hef013f);
    mcoreClass.set_mregs(32'h135, 32'h0);
    mcoreClass.set_mregs(32'h136, 32'h0);
    mcoreClass.set_mregs(32'h137, 32'h0);
    mcoreClass.set_mregs(32'h138, 32'h201000);
    mcoreClass.set_mregs(32'h139, 32'h0);
    mcoreClass.set_mregs(32'h13a, 32'h0);
    mcoreClass.set_mregs(32'h13b, 32'h0);
    mcoreClass.set_mregs(32'h13c, 32'h201000);
    mcoreClass.set_mregs(32'h13d, 32'h0);
    mcoreClass.set_mregs(32'h13e, 32'h0);
    mcoreClass.set_mregs(32'h13f, 32'h0);
    mcoreClass.set_mregs(32'h140, 32'h0);
    mcoreClass.set_mregs(32'h141, 32'h0);
    mcoreClass.set_mregs(32'h142, 32'h0);
    mcoreClass.set_mregs(32'h143, 32'h0);
    mcoreClass.set_mregs(32'h144, 32'h0);
    mcoreClass.set_mregs(32'h145, 32'h0);
    mcoreClass.set_mregs(32'h146, 32'h0);
    mcoreClass.set_mregs(32'h147, 32'h0);
    mcoreClass.set_mregs(32'h148, 32'h0);
    mcoreClass.set_mregs(32'h149, 32'h0);
    mcoreClass.set_mregs(32'h14a, 32'h0);
    mcoreClass.set_mregs(32'h14b, 32'h0);
    mcoreClass.set_mregs(32'h14c, 32'h0);
    mcoreClass.set_mregs(32'h14d, 32'h0);
    mcoreClass.set_mregs(32'h14e, 32'h0);
    mcoreClass.set_mregs(32'h14f, 32'h0);
    mcoreClass.set_mregs(32'h150, 32'h0);
    mcoreClass.set_mregs(32'h151, 32'h0);
    mcoreClass.set_mregs(32'h152, 32'h0);
    mcoreClass.set_mregs(32'h153, 32'h0);
    mcoreClass.set_mregs(32'h154, 32'h0);
    mcoreClass.set_mregs(32'h155, 32'h0);
    mcoreClass.set_mregs(32'h156, 32'h0);
    mcoreClass.set_mregs(32'h157, 32'h0);
    mcoreClass.set_mregs(32'h158, 32'h0);
    mcoreClass.set_mregs(32'h159, 32'h0);
    mcoreClass.set_mregs(32'h15a, 32'h0);
    mcoreClass.set_mregs(32'h15b, 32'h0);
    mcoreClass.set_mregs(32'h15c, 32'h0);
    mcoreClass.set_mregs(32'h15d, 32'h0);
    mcoreClass.set_mregs(32'h15e, 32'h0);
    mcoreClass.set_mregs(32'h15f, 32'h0);
    mcoreClass.set_mregs(32'h160, 32'h0);
    mcoreClass.set_mregs(32'h161, 32'h0);
    mcoreClass.set_mregs(32'h162, 32'h0);
    mcoreClass.set_mregs(32'h163, 32'h0);
    mcoreClass.set_mregs(32'h164, 32'h0);
    mcoreClass.set_mregs(32'h165, 32'h0);
    mcoreClass.set_mregs(32'h166, 32'h0);
    mcoreClass.set_mregs(32'h167, 32'h0);
    mcoreClass.set_mregs(32'h168, 32'h0);
    mcoreClass.set_mregs(32'h169, 32'h0);
    mcoreClass.set_mregs(32'h16a, 32'h0);
    mcoreClass.set_mregs(32'h16b, 32'h0);
    mcoreClass.set_mregs(32'h16c, 32'h0);
    mcoreClass.set_mregs(32'h16d, 32'h0);
    mcoreClass.set_mregs(32'h16e, 32'h0);
    mcoreClass.set_mregs(32'h16f, 32'h0);
    mcoreClass.set_mregs(32'h170, 32'h0);
    mcoreClass.set_mregs(32'h171, 32'h0);
    mcoreClass.set_mregs(32'h172, 32'h0);
    mcoreClass.set_mregs(32'h173, 32'h0);
    mcoreClass.set_mregs(32'h174, 32'h0);
    mcoreClass.set_mregs(32'h175, 32'h0);
    mcoreClass.set_mregs(32'h176, 32'h0);
    mcoreClass.set_mregs(32'h177, 32'h0);
    mcoreClass.set_mregs(32'h178, 32'h0);
    mcoreClass.set_mregs(32'h179, 32'h0);
    mcoreClass.set_mregs(32'h17a, 32'h0);
    mcoreClass.set_mregs(32'h17b, 32'h0);
    mcoreClass.set_mregs(32'h17c, 32'h0);
    mcoreClass.set_mregs(32'h17d, 32'h0);
    mcoreClass.set_mregs(32'h17e, 32'h0);
    mcoreClass.set_mregs(32'h17f, 32'h0);
    mcoreClass.set_mregs(32'h180, 32'h0);
    mcoreClass.set_mregs(32'h181, 32'h0);
    mcoreClass.set_mregs(32'h182, 32'h0);
    mcoreClass.set_mregs(32'h183, 32'h0);
    mcoreClass.set_mregs(32'h184, 32'h0);
    mcoreClass.set_mregs(32'h185, 32'h0);
    mcoreClass.set_mregs(32'h186, 32'h0);
    mcoreClass.set_mregs(32'h187, 32'h0);
    mcoreClass.set_mregs(32'h188, 32'h0);
    mcoreClass.set_mregs(32'h189, 32'h0);
    mcoreClass.set_mregs(32'h18a, 32'h0);
    mcoreClass.set_mregs(32'h18b, 32'h0);
    mcoreClass.set_mregs(32'h18c, 32'h0);
    mcoreClass.set_mregs(32'h18d, 32'h0);
    mcoreClass.set_mregs(32'h18e, 32'h0);
    mcoreClass.set_mregs(32'h18f, 32'h0);
    mcoreClass.set_mregs(32'h190, 32'h0);
    mcoreClass.set_mregs(32'h191, 32'h0);
    mcoreClass.set_mregs(32'h192, 32'h0);
    mcoreClass.set_mregs(32'h193, 32'h0);
    mcoreClass.set_mregs(32'h194, 32'h0);
    mcoreClass.set_mregs(32'h195, 32'h0);
    mcoreClass.set_mregs(32'h196, 32'h0);
    mcoreClass.set_mregs(32'h197, 32'h0);
    mcoreClass.set_mregs(32'h198, 32'h0);
    mcoreClass.set_mregs(32'h199, 32'h0);
    mcoreClass.set_mregs(32'h19a, 32'h0);
    mcoreClass.set_mregs(32'h19b, 32'h0);
    mcoreClass.set_mregs(32'h19c, 32'h0);
    mcoreClass.set_mregs(32'h19d, 32'h0);
    mcoreClass.set_mregs(32'h19e, 32'h0);
    mcoreClass.set_mregs(32'h19f, 32'h0);
    mcoreClass.set_mregs(32'h1a0, 32'h0);
    mcoreClass.set_mregs(32'h1a1, 32'h0);
    mcoreClass.set_mregs(32'h1a2, 32'h0);
    mcoreClass.set_mregs(32'h1a3, 32'h0);
    mcoreClass.set_mregs(32'h1a4, 32'h0);
    mcoreClass.set_mregs(32'h1a5, 32'h0);
    mcoreClass.set_mregs(32'h1a6, 32'h0);
    mcoreClass.set_mregs(32'h1a7, 32'h0);
    mcoreClass.set_mregs(32'h1a8, 32'h0);
    mcoreClass.set_mregs(32'h1a9, 32'h0);
    mcoreClass.set_mregs(32'h1aa, 32'h0);
    mcoreClass.set_mregs(32'h1ab, 32'h0);
    mcoreClass.set_mregs(32'h1ac, 32'h0);
    mcoreClass.set_mregs(32'h1ad, 32'h0);
    mcoreClass.set_mregs(32'h1ae, 32'h0);
    mcoreClass.set_mregs(32'h1af, 32'h0);
    mcoreClass.set_mregs(32'h1b0, 32'h0);
    mcoreClass.set_mregs(32'h1b1, 32'h0);
    mcoreClass.set_mregs(32'h1b2, 32'h0);
    mcoreClass.set_mregs(32'h1b3, 32'h0);
    mcoreClass.set_mregs(32'h1b4, 32'h0);
    mcoreClass.set_mregs(32'h1b5, 32'h0);
    mcoreClass.set_mregs(32'h1b6, 32'h0);
    mcoreClass.set_mregs(32'h1b7, 32'h0);
    mcoreClass.set_mregs(32'h1b8, 32'h0);
    mcoreClass.set_mregs(32'h1b9, 32'h0);
    mcoreClass.set_mregs(32'h1ba, 32'h0);
    mcoreClass.set_mregs(32'h1bb, 32'h0);
    mcoreClass.set_mregs(32'h1bc, 32'h0);
    mcoreClass.set_mregs(32'h1bd, 32'h0);
    mcoreClass.set_mregs(32'h1be, 32'h0);
    mcoreClass.set_mregs(32'h1bf, 32'h0);
    mcoreClass.set_mregs(32'h1c0, 32'h0);
    mcoreClass.set_mregs(32'h1c1, 32'h0);
    mcoreClass.set_mregs(32'h1c2, 32'h0);
    mcoreClass.set_mregs(32'h1c3, 32'h0);
    mcoreClass.set_mregs(32'h1c4, 32'h0);
    mcoreClass.set_mregs(32'h1c5, 32'h0);
    mcoreClass.set_mregs(32'h1c6, 32'h0);
    mcoreClass.set_mregs(32'h1c7, 32'h0);
    mcoreClass.set_mregs(32'h1c8, 32'h0);
    mcoreClass.set_mregs(32'h1c9, 32'h0);
    mcoreClass.set_mregs(32'h1ca, 32'h0);
    mcoreClass.set_mregs(32'h1cb, 32'h0);
    mcoreClass.set_mregs(32'h1cc, 32'h0);
    mcoreClass.set_mregs(32'h1cd, 32'h0);
    mcoreClass.set_mregs(32'h1ce, 32'h0);
    mcoreClass.set_mregs(32'h1cf, 32'h0);
    mcoreClass.set_mregs(32'h1d0, 32'h0);
    mcoreClass.set_mregs(32'h1d1, 32'h0);
    mcoreClass.set_mregs(32'h1d2, 32'h0);
    mcoreClass.set_mregs(32'h1d3, 32'h0);
    mcoreClass.set_mregs(32'h1d4, 32'h0);
    mcoreClass.set_mregs(32'h1d5, 32'h0);
    mcoreClass.set_mregs(32'h1d6, 32'h0);
    mcoreClass.set_mregs(32'h1d7, 32'h0);
    mcoreClass.set_mregs(32'h1d8, 32'h0);
    mcoreClass.set_mregs(32'h1d9, 32'h0);
    mcoreClass.set_mregs(32'h1da, 32'h0);
    mcoreClass.set_mregs(32'h1db, 32'h0);
    mcoreClass.set_mregs(32'h1dc, 32'h0);
    mcoreClass.set_mregs(32'h1dd, 32'h0);
    mcoreClass.set_mregs(32'h1de, 32'h0);
    mcoreClass.set_mregs(32'h1df, 32'h0);
    mcoreClass.set_mregs(32'h1e0, 32'h0);
    mcoreClass.set_mregs(32'h1e1, 32'h0);
    mcoreClass.set_mregs(32'h1e2, 32'h0);
    mcoreClass.set_mregs(32'h1e3, 32'h0);
    mcoreClass.set_mregs(32'h1e4, 32'h0);
    mcoreClass.set_mregs(32'h1e5, 32'h0);
    mcoreClass.set_mregs(32'h1e6, 32'h0);
    mcoreClass.set_mregs(32'h1e7, 32'h0);
    mcoreClass.set_mregs(32'h1e8, 32'h0);
    mcoreClass.set_mregs(32'h1e9, 32'h0);
    mcoreClass.set_mregs(32'h1ea, 32'h0);
    mcoreClass.set_mregs(32'h1eb, 32'h0);
    mcoreClass.set_mregs(32'h1ec, 32'h0);
    mcoreClass.set_mregs(32'h1ed, 32'h0);
    mcoreClass.set_mregs(32'h1ee, 32'h0);
    mcoreClass.set_mregs(32'h1ef, 32'h0);
    mcoreClass.set_mregs(32'h1f0, 32'h0);
    mcoreClass.set_mregs(32'h1f1, 32'h0);
    mcoreClass.set_mregs(32'h1f2, 32'h0);
    mcoreClass.set_mregs(32'h1f3, 32'h0);
    mcoreClass.set_mregs(32'h1f4, 32'h0);
    mcoreClass.set_mregs(32'h1f5, 32'h0);
    mcoreClass.set_mregs(32'h1f6, 32'h0);
    mcoreClass.set_mregs(32'h1f7, 32'h0);
    mcoreClass.set_mregs(32'h1f8, 32'h0);
    mcoreClass.set_mregs(32'h1f9, 32'h0);
    mcoreClass.set_mregs(32'h1fa, 32'h0);
    mcoreClass.set_mregs(32'h1fb, 32'h0);
    mcoreClass.set_mregs(32'h1fc, 32'h0);
    mcoreClass.set_mregs(32'h1fd, 32'h0);
    mcoreClass.set_mregs(32'h1fe, 32'h0);
    mcoreClass.set_mregs(32'h1ff, 32'h0);
    mcoreClass.set_mregs(32'h200, 32'h0);
    mcoreClass.set_mregs(32'h201, 32'h0);
    mcoreClass.set_mregs(32'h202, 32'h0);
    mcoreClass.set_mregs(32'h203, 32'h0);
    mcoreClass.set_mregs(32'h204, 32'h0);
    mcoreClass.set_mregs(32'h205, 32'h0);
    mcoreClass.set_mregs(32'h206, 32'h0);
    mcoreClass.set_mregs(32'h207, 32'h0);
    mcoreClass.set_mregs(32'h208, 32'h0);
    mcoreClass.set_mregs(32'h209, 32'h0);
    mcoreClass.set_mregs(32'h20a, 32'h0);
    mcoreClass.set_mregs(32'h20b, 32'h0);
    mcoreClass.set_mregs(32'h20c, 32'h0);
    mcoreClass.set_mregs(32'h20d, 32'h0);
    mcoreClass.set_mregs(32'h20e, 32'h0);
    mcoreClass.set_mregs(32'h20f, 32'h0);
    mcoreClass.set_mregs(32'h210, 32'h0);
    mcoreClass.set_mregs(32'h211, 32'h0);
    mcoreClass.set_mregs(32'h212, 32'h0);
    mcoreClass.set_mregs(32'h213, 32'h0);
    mcoreClass.set_mregs(32'h214, 32'h0);
    mcoreClass.set_mregs(32'h215, 32'h0);
    mcoreClass.set_mregs(32'h216, 32'h0);
    mcoreClass.set_mregs(32'h217, 32'h0);
    mcoreClass.set_mregs(32'h218, 32'hffff8000);
    mcoreClass.set_mregs(32'h219, 32'h0);
    mcoreClass.set_mregs(32'h21a, 32'h0);
    mcoreClass.set_mregs(32'h21b, 32'h0);
    mcoreClass.set_mregs(32'h21c, 32'hfffffff);
    mcoreClass.set_mregs(32'h21d, 32'h0);
    mcoreClass.set_mregs(32'h21e, 32'h0);
    mcoreClass.set_mregs(32'h21f, 32'h0);
    mcoreClass.set_mregs(32'h220, 32'h0);
    mcoreClass.set_mregs(32'h221, 32'h0);
    mcoreClass.set_mregs(32'h222, 32'h0);
    mcoreClass.set_mregs(32'h223, 32'h0);
    mcoreClass.set_mregs(32'h224, 32'h0);
    mcoreClass.set_mregs(32'h225, 32'h0);
    mcoreClass.set_mregs(32'h226, 32'h0);
    mcoreClass.set_mregs(32'h227, 32'h0);
    mcoreClass.set_mregs(32'h228, 32'h0);
    mcoreClass.set_mregs(32'h229, 32'h0);
    mcoreClass.set_mregs(32'h22a, 32'h0);
    mcoreClass.set_mregs(32'h22b, 32'h0);
    mcoreClass.set_mregs(32'h22c, 32'h0);
    mcoreClass.set_mregs(32'h22d, 32'h0);
    mcoreClass.set_mregs(32'h22e, 32'h0);
    mcoreClass.set_mregs(32'h22f, 32'h0);
    mcoreClass.set_mregs(32'h230, 32'h0);
    mcoreClass.set_mregs(32'h231, 32'h0);
    mcoreClass.set_mregs(32'h232, 32'h0);
    mcoreClass.set_mregs(32'h233, 32'h0);
    mcoreClass.set_mregs(32'h234, 32'h0);
    mcoreClass.set_mregs(32'h235, 32'h0);
    mcoreClass.set_mregs(32'h236, 32'h0);
    mcoreClass.set_mregs(32'h237, 32'h0);
    mcoreClass.set_mregs(32'h238, 32'hffffffff);
    mcoreClass.set_mregs(32'h239, 32'h0);
    mcoreClass.set_mregs(32'h23a, 32'h0);
    mcoreClass.set_mregs(32'h23b, 32'h0);
    mcoreClass.set_mregs(32'h23c, 32'h7fffffff);
    mcoreClass.set_mregs(32'h23d, 32'h0);
    mcoreClass.set_mregs(32'h23e, 32'hfffffffc);
    mcoreClass.set_mregs(32'h23f, 32'h0);
    mcoreClass.set_mregs(32'h240, 32'h0);
    mcoreClass.set_mregs(32'h241, 32'h0);
    mcoreClass.set_mregs(32'h242, 32'h0);
    mcoreClass.set_mregs(32'h243, 32'h0);
    mcoreClass.set_mregs(32'h244, 32'h0);
    mcoreClass.set_mregs(32'h245, 32'h0);
    mcoreClass.set_mregs(32'h246, 32'h0);
    mcoreClass.set_mregs(32'h247, 32'h0);
    mcoreClass.set_mregs(32'h248, 32'h0);
    mcoreClass.set_mregs(32'h249, 32'h0);
    mcoreClass.set_mregs(32'h24a, 32'h0);
    mcoreClass.set_mregs(32'h24b, 32'h0);
    mcoreClass.set_mregs(32'h24c, 32'h0);
    mcoreClass.set_mregs(32'h24d, 32'h0);
    mcoreClass.set_mregs(32'h24e, 32'h0);
    mcoreClass.set_mregs(32'h24f, 32'h0);
    mcoreClass.set_mregs(32'h250, 32'h0);
    mcoreClass.set_mregs(32'h251, 32'h0);
    mcoreClass.set_mregs(32'h252, 32'h0);
    mcoreClass.set_mregs(32'h253, 32'h0);
    mcoreClass.set_mregs(32'h254, 32'h0);
    mcoreClass.set_mregs(32'h255, 32'h0);
    mcoreClass.set_mregs(32'h256, 32'h0);
    mcoreClass.set_mregs(32'h257, 32'h0);
    mcoreClass.set_mregs(32'h258, 32'h0);
    mcoreClass.set_mregs(32'h259, 32'h0);
    mcoreClass.set_mregs(32'h25a, 32'h0);
    mcoreClass.set_mregs(32'h25b, 32'h0);
    mcoreClass.set_mregs(32'h25c, 32'h0);
    mcoreClass.set_mregs(32'h25d, 32'h0);
    mcoreClass.set_mregs(32'h25e, 32'h0);
    mcoreClass.set_mregs(32'h25f, 32'h0);
    mcoreClass.set_mregs(32'h260, 32'h0);
    mcoreClass.set_mregs(32'h261, 32'h0);
    mcoreClass.set_mregs(32'h262, 32'h0);
    mcoreClass.set_mregs(32'h263, 32'h0);
    mcoreClass.set_mregs(32'h264, 32'h0);
    mcoreClass.set_mregs(32'h265, 32'h0);
    mcoreClass.set_mregs(32'h266, 32'h0);
    mcoreClass.set_mregs(32'h267, 32'h0);
    mcoreClass.set_mregs(32'h268, 32'h0);
    mcoreClass.set_mregs(32'h269, 32'h0);
    mcoreClass.set_mregs(32'h26a, 32'h0);
    mcoreClass.set_mregs(32'h26b, 32'h0);
    mcoreClass.set_mregs(32'h26c, 32'h0);
    mcoreClass.set_mregs(32'h26d, 32'h0);
    mcoreClass.set_mregs(32'h26e, 32'h0);
    mcoreClass.set_mregs(32'h26f, 32'h0);
    mcoreClass.set_mregs(32'h270, 32'h0);
    mcoreClass.set_mregs(32'h271, 32'h0);
    mcoreClass.set_mregs(32'h272, 32'h0);
    mcoreClass.set_mregs(32'h273, 32'h0);
    mcoreClass.set_mregs(32'h274, 32'h0);
    mcoreClass.set_mregs(32'h275, 32'h0);
    mcoreClass.set_mregs(32'h276, 32'h0);
    mcoreClass.set_mregs(32'h277, 32'h0);
    mcoreClass.set_mregs(32'h278, 32'h0);
    mcoreClass.set_mregs(32'h279, 32'h0);
    mcoreClass.set_mregs(32'h27a, 32'h0);
    mcoreClass.set_mregs(32'h27b, 32'h0);
    mcoreClass.set_mregs(32'h27c, 32'h0);
    mcoreClass.set_mregs(32'h27d, 32'h0);
    mcoreClass.set_mregs(32'h27e, 32'h0);
    mcoreClass.set_mregs(32'h27f, 32'h0);
    mcoreClass.set_mregs(32'h280, 32'h0);
    mcoreClass.set_mregs(32'h281, 32'h0);
    mcoreClass.set_mregs(32'h282, 32'h0);
    mcoreClass.set_mregs(32'h283, 32'h0);
    mcoreClass.set_mregs(32'h284, 32'h0);
    mcoreClass.set_mregs(32'h285, 32'h0);
    mcoreClass.set_mregs(32'h286, 32'h0);
    mcoreClass.set_mregs(32'h287, 32'h0);
    mcoreClass.set_mregs(32'h288, 32'h0);
    mcoreClass.set_mregs(32'h289, 32'h0);
    mcoreClass.set_mregs(32'h28a, 32'h0);
    mcoreClass.set_mregs(32'h28b, 32'h0);
    mcoreClass.set_mregs(32'h28c, 32'h0);
    mcoreClass.set_mregs(32'h28d, 32'h0);
    mcoreClass.set_mregs(32'h28e, 32'h0);
    mcoreClass.set_mregs(32'h28f, 32'h0);
    mcoreClass.set_mregs(32'h290, 32'h0);
    mcoreClass.set_mregs(32'h291, 32'h0);
    mcoreClass.set_mregs(32'h292, 32'h0);
    mcoreClass.set_mregs(32'h293, 32'h0);
    mcoreClass.set_mregs(32'h294, 32'h0);
    mcoreClass.set_mregs(32'h295, 32'h0);
    mcoreClass.set_mregs(32'h296, 32'h0);
    mcoreClass.set_mregs(32'h297, 32'h0);
    mcoreClass.set_mregs(32'h298, 32'h0);
    mcoreClass.set_mregs(32'h299, 32'h0);
    mcoreClass.set_mregs(32'h29a, 32'h0);
    mcoreClass.set_mregs(32'h29b, 32'h0);
    mcoreClass.set_mregs(32'h29c, 32'h0);
    mcoreClass.set_mregs(32'h29d, 32'h0);
    mcoreClass.set_mregs(32'h29e, 32'h0);
    mcoreClass.set_mregs(32'h29f, 32'h0);
    mcoreClass.set_mregs(32'h2a0, 32'h0);
    mcoreClass.set_mregs(32'h2a1, 32'h0);
    mcoreClass.set_mregs(32'h2a2, 32'h0);
    mcoreClass.set_mregs(32'h2a3, 32'h0);
    mcoreClass.set_mregs(32'h2a4, 32'h0);
    mcoreClass.set_mregs(32'h2a5, 32'h0);
    mcoreClass.set_mregs(32'h2a6, 32'h0);
    mcoreClass.set_mregs(32'h2a7, 32'h0);
    mcoreClass.set_mregs(32'h2a8, 32'h0);
    mcoreClass.set_mregs(32'h2a9, 32'h0);
    mcoreClass.set_mregs(32'h2aa, 32'h0);
    mcoreClass.set_mregs(32'h2ab, 32'h0);
    mcoreClass.set_mregs(32'h2ac, 32'h0);
    mcoreClass.set_mregs(32'h2ad, 32'h0);
    mcoreClass.set_mregs(32'h2ae, 32'h0);
    mcoreClass.set_mregs(32'h2af, 32'h0);
    mcoreClass.set_mregs(32'h2b0, 32'h0);
    mcoreClass.set_mregs(32'h2b1, 32'h0);
    mcoreClass.set_mregs(32'h2b2, 32'h0);
    mcoreClass.set_mregs(32'h2b3, 32'h0);
    mcoreClass.set_mregs(32'h2b4, 32'h0);
    mcoreClass.set_mregs(32'h2b5, 32'h0);
    mcoreClass.set_mregs(32'h2b6, 32'h0);
    mcoreClass.set_mregs(32'h2b7, 32'h0);
    mcoreClass.set_mregs(32'h2b8, 32'h0);
    mcoreClass.set_mregs(32'h2b9, 32'h0);
    mcoreClass.set_mregs(32'h2ba, 32'h0);
    mcoreClass.set_mregs(32'h2bb, 32'h0);
    mcoreClass.set_mregs(32'h2bc, 32'h0);
    mcoreClass.set_mregs(32'h2bd, 32'h0);
    mcoreClass.set_mregs(32'h2be, 32'h0);
    mcoreClass.set_mregs(32'h2bf, 32'h0);
    mcoreClass.set_mregs(32'h2c0, 32'h0);
    mcoreClass.set_mregs(32'h2c1, 32'h0);
    mcoreClass.set_mregs(32'h2c2, 32'h0);
    mcoreClass.set_mregs(32'h2c3, 32'h0);
    mcoreClass.set_mregs(32'h2c4, 32'h0);
    mcoreClass.set_mregs(32'h2c5, 32'h0);
    mcoreClass.set_mregs(32'h2c6, 32'h0);
    mcoreClass.set_mregs(32'h2c7, 32'h0);
    mcoreClass.set_mregs(32'h2c8, 32'h0);
    mcoreClass.set_mregs(32'h2c9, 32'h0);
    mcoreClass.set_mregs(32'h2ca, 32'h0);
    mcoreClass.set_mregs(32'h2cb, 32'h0);
    mcoreClass.set_mregs(32'h2cc, 32'h0);
    mcoreClass.set_mregs(32'h2cd, 32'h0);
    mcoreClass.set_mregs(32'h2ce, 32'h0);
    mcoreClass.set_mregs(32'h2cf, 32'h0);
    mcoreClass.set_mregs(32'h2d0, 32'h0);
    mcoreClass.set_mregs(32'h2d1, 32'h0);
    mcoreClass.set_mregs(32'h2d2, 32'h0);
    mcoreClass.set_mregs(32'h2d3, 32'h0);
    mcoreClass.set_mregs(32'h2d4, 32'h0);
    mcoreClass.set_mregs(32'h2d5, 32'h0);
    mcoreClass.set_mregs(32'h2d6, 32'h0);
    mcoreClass.set_mregs(32'h2d7, 32'h0);
    mcoreClass.set_mregs(32'h2d8, 32'h0);
    mcoreClass.set_mregs(32'h2d9, 32'h0);
    mcoreClass.set_mregs(32'h2da, 32'h0);
    mcoreClass.set_mregs(32'h2db, 32'h0);
    mcoreClass.set_mregs(32'h2dc, 32'h0);
    mcoreClass.set_mregs(32'h2dd, 32'h0);
    mcoreClass.set_mregs(32'h2de, 32'h0);
    mcoreClass.set_mregs(32'h2df, 32'h0);
    mcoreClass.set_mregs(32'h2e0, 32'h0);
    mcoreClass.set_mregs(32'h2e1, 32'h0);
    mcoreClass.set_mregs(32'h2e2, 32'h0);
    mcoreClass.set_mregs(32'h2e3, 32'h0);
    mcoreClass.set_mregs(32'h2e4, 32'h0);
    mcoreClass.set_mregs(32'h2e5, 32'h0);
    mcoreClass.set_mregs(32'h2e6, 32'h0);
    mcoreClass.set_mregs(32'h2e7, 32'h0);
    mcoreClass.set_mregs(32'h2e8, 32'h0);
    mcoreClass.set_mregs(32'h2e9, 32'h0);
    mcoreClass.set_mregs(32'h2ea, 32'h0);
    mcoreClass.set_mregs(32'h2eb, 32'h0);
    mcoreClass.set_mregs(32'h2ec, 32'h0);
    mcoreClass.set_mregs(32'h2ed, 32'h0);
    mcoreClass.set_mregs(32'h2ee, 32'h0);
    mcoreClass.set_mregs(32'h2ef, 32'h0);
    mcoreClass.set_mregs(32'h2f0, 32'h0);
    mcoreClass.set_mregs(32'h2f1, 32'h0);
    mcoreClass.set_mregs(32'h2f2, 32'h0);
    mcoreClass.set_mregs(32'h2f3, 32'h0);
    mcoreClass.set_mregs(32'h2f4, 32'h0);
    mcoreClass.set_mregs(32'h2f5, 32'h0);
    mcoreClass.set_mregs(32'h2f6, 32'h0);
    mcoreClass.set_mregs(32'h2f7, 32'h0);
    mcoreClass.set_mregs(32'h2f8, 32'h0);
    mcoreClass.set_mregs(32'h2f9, 32'h0);
    mcoreClass.set_mregs(32'h2fa, 32'h0);
    mcoreClass.set_mregs(32'h2fb, 32'h0);
    mcoreClass.set_mregs(32'h2fc, 32'h0);
    mcoreClass.set_mregs(32'h2fd, 32'h0);
    mcoreClass.set_mregs(32'h2fe, 32'h0);
    mcoreClass.set_mregs(32'h2ff, 32'h0);
    mcoreClass.set_mregs(32'h300, 32'h0);
    mcoreClass.set_mregs(32'h301, 32'h0);
    mcoreClass.set_mregs(32'h302, 32'h0);
    mcoreClass.set_mregs(32'h303, 32'h0);
    mcoreClass.set_mregs(32'h304, 32'h0);
    mcoreClass.set_mregs(32'h305, 32'h0);
    mcoreClass.set_mregs(32'h306, 32'h0);
    mcoreClass.set_mregs(32'h307, 32'h0);
    mcoreClass.set_mregs(32'h308, 32'h0);
    mcoreClass.set_mregs(32'h309, 32'h0);
    mcoreClass.set_mregs(32'h30a, 32'h0);
    mcoreClass.set_mregs(32'h30b, 32'h0);
    mcoreClass.set_mregs(32'h30c, 32'h0);
    mcoreClass.set_mregs(32'h30d, 32'h0);
    mcoreClass.set_mregs(32'h30e, 32'h0);
    mcoreClass.set_mregs(32'h30f, 32'h0);
    mcoreClass.set_mregs(32'h310, 32'h0);
    mcoreClass.set_mregs(32'h311, 32'h0);
    mcoreClass.set_mregs(32'h312, 32'h0);
    mcoreClass.set_mregs(32'h313, 32'h0);
    mcoreClass.set_mregs(32'h314, 32'h0);
    mcoreClass.set_mregs(32'h315, 32'h0);
    mcoreClass.set_mregs(32'h316, 32'h0);
    mcoreClass.set_mregs(32'h317, 32'h0);
    mcoreClass.set_mregs(32'h318, 32'h0);
    mcoreClass.set_mregs(32'h319, 32'h0);
    mcoreClass.set_mregs(32'h31a, 32'h0);
    mcoreClass.set_mregs(32'h31b, 32'h0);
    mcoreClass.set_mregs(32'h31c, 32'h0);
    mcoreClass.set_mregs(32'h31d, 32'h0);
    mcoreClass.set_mregs(32'h31e, 32'h0);
    mcoreClass.set_mregs(32'h31f, 32'h0);
    mcoreClass.set_mregs(32'h320, 32'h0);
    mcoreClass.set_mregs(32'h321, 32'h0);
    mcoreClass.set_mregs(32'h322, 32'h0);
    mcoreClass.set_mregs(32'h323, 32'h0);
    mcoreClass.set_mregs(32'h324, 32'h0);
    mcoreClass.set_mregs(32'h325, 32'h0);
    mcoreClass.set_mregs(32'h326, 32'h0);
    mcoreClass.set_mregs(32'h327, 32'h0);
    mcoreClass.set_mregs(32'h328, 32'h0);
    mcoreClass.set_mregs(32'h329, 32'h0);
    mcoreClass.set_mregs(32'h32a, 32'h0);
    mcoreClass.set_mregs(32'h32b, 32'h0);
    mcoreClass.set_mregs(32'h32c, 32'h0);
    mcoreClass.set_mregs(32'h32d, 32'h0);
    mcoreClass.set_mregs(32'h32e, 32'h0);
    mcoreClass.set_mregs(32'h32f, 32'h0);
    mcoreClass.set_mregs(32'h330, 32'h0);
    mcoreClass.set_mregs(32'h331, 32'h0);
    mcoreClass.set_mregs(32'h332, 32'h0);
    mcoreClass.set_mregs(32'h333, 32'h0);
    mcoreClass.set_mregs(32'h334, 32'h0);
    mcoreClass.set_mregs(32'h335, 32'h0);
    mcoreClass.set_mregs(32'h336, 32'h0);
    mcoreClass.set_mregs(32'h337, 32'h0);
    mcoreClass.set_mregs(32'h338, 32'h0);
    mcoreClass.set_mregs(32'h339, 32'h0);
    mcoreClass.set_mregs(32'h33a, 32'h0);
    mcoreClass.set_mregs(32'h33b, 32'h0);
    mcoreClass.set_mregs(32'h33c, 32'h0);
    mcoreClass.set_mregs(32'h33d, 32'h0);
    mcoreClass.set_mregs(32'h33e, 32'h0);
    mcoreClass.set_mregs(32'h33f, 32'h0);
    mcoreClass.set_mregs(32'h340, 32'h0);
    mcoreClass.set_mregs(32'h341, 32'h0);
    mcoreClass.set_mregs(32'h342, 32'h0);
    mcoreClass.set_mregs(32'h343, 32'h0);
    mcoreClass.set_mregs(32'h344, 32'h0);
    mcoreClass.set_mregs(32'h345, 32'h0);
    mcoreClass.set_mregs(32'h346, 32'h0);
    mcoreClass.set_mregs(32'h347, 32'h0);
    mcoreClass.set_mregs(32'h348, 32'h0);
    mcoreClass.set_mregs(32'h349, 32'h0);
    mcoreClass.set_mregs(32'h34a, 32'h0);
    mcoreClass.set_mregs(32'h34b, 32'h0);
    mcoreClass.set_mregs(32'h34c, 32'h0);
    mcoreClass.set_mregs(32'h34d, 32'h0);
    mcoreClass.set_mregs(32'h34e, 32'h0);
    mcoreClass.set_mregs(32'h34f, 32'h0);
    mcoreClass.set_mregs(32'h350, 32'h0);
    mcoreClass.set_mregs(32'h351, 32'h0);
    mcoreClass.set_mregs(32'h352, 32'h0);
    mcoreClass.set_mregs(32'h353, 32'h0);
    mcoreClass.set_mregs(32'h354, 32'h0);
    mcoreClass.set_mregs(32'h355, 32'h0);
    mcoreClass.set_mregs(32'h356, 32'h0);
    mcoreClass.set_mregs(32'h357, 32'h0);
    mcoreClass.set_mregs(32'h358, 32'h0);
    mcoreClass.set_mregs(32'h359, 32'h0);
    mcoreClass.set_mregs(32'h35a, 32'h0);
    mcoreClass.set_mregs(32'h35b, 32'h0);
    mcoreClass.set_mregs(32'h35c, 32'h0);
    mcoreClass.set_mregs(32'h35d, 32'h0);
    mcoreClass.set_mregs(32'h35e, 32'h0);
    mcoreClass.set_mregs(32'h35f, 32'h0);
    mcoreClass.set_mregs(32'h360, 32'h0);
    mcoreClass.set_mregs(32'h361, 32'h0);
    mcoreClass.set_mregs(32'h362, 32'h0);
    mcoreClass.set_mregs(32'h363, 32'h0);
    mcoreClass.set_mregs(32'h364, 32'h0);
    mcoreClass.set_mregs(32'h365, 32'h0);
    mcoreClass.set_mregs(32'h366, 32'h0);
    mcoreClass.set_mregs(32'h367, 32'h0);
    mcoreClass.set_mregs(32'h368, 32'h0);
    mcoreClass.set_mregs(32'h369, 32'h0);
    mcoreClass.set_mregs(32'h36a, 32'h0);
    mcoreClass.set_mregs(32'h36b, 32'h0);
    mcoreClass.set_mregs(32'h36c, 32'h0);
    mcoreClass.set_mregs(32'h36d, 32'h0);
    mcoreClass.set_mregs(32'h36e, 32'h0);
    mcoreClass.set_mregs(32'h36f, 32'h0);
    mcoreClass.set_mregs(32'h370, 32'h0);
    mcoreClass.set_mregs(32'h371, 32'h0);
    mcoreClass.set_mregs(32'h372, 32'h0);
    mcoreClass.set_mregs(32'h373, 32'h0);
    mcoreClass.set_mregs(32'h374, 32'h0);
    mcoreClass.set_mregs(32'h375, 32'h0);
    mcoreClass.set_mregs(32'h376, 32'h0);
    mcoreClass.set_mregs(32'h377, 32'h0);
    mcoreClass.set_mregs(32'h378, 32'h0);
    mcoreClass.set_mregs(32'h379, 32'h0);
    mcoreClass.set_mregs(32'h37a, 32'h0);
    mcoreClass.set_mregs(32'h37b, 32'h0);
    mcoreClass.set_mregs(32'h37c, 32'h0);
    mcoreClass.set_mregs(32'h37d, 32'h0);
    mcoreClass.set_mregs(32'h37e, 32'h0);
    mcoreClass.set_mregs(32'h37f, 32'h0);
    mcoreClass.set_mregs(32'h380, 32'h0);
    mcoreClass.set_mregs(32'h381, 32'h0);
    mcoreClass.set_mregs(32'h382, 32'h0);
    mcoreClass.set_mregs(32'h383, 32'h0);
    mcoreClass.set_mregs(32'h384, 32'h0);
    mcoreClass.set_mregs(32'h385, 32'h0);
    mcoreClass.set_mregs(32'h386, 32'h0);
    mcoreClass.set_mregs(32'h387, 32'h0);
    mcoreClass.set_mregs(32'h388, 32'h0);
    mcoreClass.set_mregs(32'h389, 32'h0);
    mcoreClass.set_mregs(32'h38a, 32'h0);
    mcoreClass.set_mregs(32'h38b, 32'h0);
    mcoreClass.set_mregs(32'h38c, 32'h0);
    mcoreClass.set_mregs(32'h38d, 32'h0);
    mcoreClass.set_mregs(32'h38e, 32'h0);
    mcoreClass.set_mregs(32'h38f, 32'h0);
    mcoreClass.set_mregs(32'h390, 32'h0);
    mcoreClass.set_mregs(32'h391, 32'h0);
    mcoreClass.set_mregs(32'h392, 32'h0);
    mcoreClass.set_mregs(32'h393, 32'h0);
    mcoreClass.set_mregs(32'h394, 32'h0);
    mcoreClass.set_mregs(32'h395, 32'h0);
    mcoreClass.set_mregs(32'h396, 32'h0);
    mcoreClass.set_mregs(32'h397, 32'h0);
    mcoreClass.set_mregs(32'h398, 32'h0);
    mcoreClass.set_mregs(32'h399, 32'h0);
    mcoreClass.set_mregs(32'h39a, 32'h0);
    mcoreClass.set_mregs(32'h39b, 32'h0);
    mcoreClass.set_mregs(32'h39c, 32'h0);
    mcoreClass.set_mregs(32'h39d, 32'h0);
    mcoreClass.set_mregs(32'h39e, 32'h0);
    mcoreClass.set_mregs(32'h39f, 32'h0);
    mcoreClass.set_mregs(32'h3a0, 32'h0);
    mcoreClass.set_mregs(32'h3a1, 32'h0);
    mcoreClass.set_mregs(32'h3a2, 32'h0);
    mcoreClass.set_mregs(32'h3a3, 32'h0);
    mcoreClass.set_mregs(32'h3a4, 32'h0);
    mcoreClass.set_mregs(32'h3a5, 32'h0);
    mcoreClass.set_mregs(32'h3a6, 32'h0);
    mcoreClass.set_mregs(32'h3a7, 32'h0);
    mcoreClass.set_mregs(32'h3a8, 32'h0);
    mcoreClass.set_mregs(32'h3a9, 32'h0);
    mcoreClass.set_mregs(32'h3aa, 32'h0);
    mcoreClass.set_mregs(32'h3ab, 32'h0);
    mcoreClass.set_mregs(32'h3ac, 32'h0);
    mcoreClass.set_mregs(32'h3ad, 32'h0);
    mcoreClass.set_mregs(32'h3ae, 32'h0);
    mcoreClass.set_mregs(32'h3af, 32'h0);
    mcoreClass.set_mregs(32'h3b0, 32'h0);
    mcoreClass.set_mregs(32'h3b1, 32'h0);
    mcoreClass.set_mregs(32'h3b2, 32'h0);
    mcoreClass.set_mregs(32'h3b3, 32'h0);
    mcoreClass.set_mregs(32'h3b4, 32'h0);
    mcoreClass.set_mregs(32'h3b5, 32'h0);
    mcoreClass.set_mregs(32'h3b6, 32'h0);
    mcoreClass.set_mregs(32'h3b7, 32'h0);
    mcoreClass.set_mregs(32'h3b8, 32'h0);
    mcoreClass.set_mregs(32'h3b9, 32'h0);
    mcoreClass.set_mregs(32'h3ba, 32'h0);
    mcoreClass.set_mregs(32'h3bb, 32'h0);
    mcoreClass.set_mregs(32'h3bc, 32'h0);
    mcoreClass.set_mregs(32'h3bd, 32'h0);
    mcoreClass.set_mregs(32'h3be, 32'h0);
    mcoreClass.set_mregs(32'h3bf, 32'h0);
    mcoreClass.set_mregs(32'h3c0, 32'h0);
    mcoreClass.set_mregs(32'h3c1, 32'h0);
    mcoreClass.set_mregs(32'h3c2, 32'h0);
    mcoreClass.set_mregs(32'h3c3, 32'h0);
    mcoreClass.set_mregs(32'h3c4, 32'h0);
    mcoreClass.set_mregs(32'h3c5, 32'h0);
    mcoreClass.set_mregs(32'h3c6, 32'h0);
    mcoreClass.set_mregs(32'h3c7, 32'h0);
    mcoreClass.set_mregs(32'h3c8, 32'h0);
    mcoreClass.set_mregs(32'h3c9, 32'h0);
    mcoreClass.set_mregs(32'h3ca, 32'h0);
    mcoreClass.set_mregs(32'h3cb, 32'h0);
    mcoreClass.set_mregs(32'h3cc, 32'h0);
    mcoreClass.set_mregs(32'h3cd, 32'h0);
    mcoreClass.set_mregs(32'h3ce, 32'h0);
    mcoreClass.set_mregs(32'h3cf, 32'h0);
    mcoreClass.set_mregs(32'h3d0, 32'h0);
    mcoreClass.set_mregs(32'h3d1, 32'h0);
    mcoreClass.set_mregs(32'h3d2, 32'h0);
    mcoreClass.set_mregs(32'h3d3, 32'h0);
    mcoreClass.set_mregs(32'h3d4, 32'h0);
    mcoreClass.set_mregs(32'h3d5, 32'h0);
    mcoreClass.set_mregs(32'h3d6, 32'h0);
    mcoreClass.set_mregs(32'h3d7, 32'h0);
    mcoreClass.set_mregs(32'h3d8, 32'h0);
    mcoreClass.set_mregs(32'h3d9, 32'h0);
    mcoreClass.set_mregs(32'h3da, 32'h0);
    mcoreClass.set_mregs(32'h3db, 32'h0);
    mcoreClass.set_mregs(32'h3dc, 32'h0);
    mcoreClass.set_mregs(32'h3dd, 32'h0);
    mcoreClass.set_mregs(32'h3de, 32'h0);
    mcoreClass.set_mregs(32'h3df, 32'h0);
    mcoreClass.set_mregs(32'h3e0, 32'h0);
    mcoreClass.set_mregs(32'h3e1, 32'h0);
    mcoreClass.set_mregs(32'h3e2, 32'h0);
    mcoreClass.set_mregs(32'h3e3, 32'h0);
    mcoreClass.set_mregs(32'h3e4, 32'h0);
    mcoreClass.set_mregs(32'h3e5, 32'h0);
    mcoreClass.set_mregs(32'h3e6, 32'h0);
    mcoreClass.set_mregs(32'h3e7, 32'h0);
    mcoreClass.set_mregs(32'h3e8, 32'h0);
    mcoreClass.set_mregs(32'h3e9, 32'h0);
    mcoreClass.set_mregs(32'h3ea, 32'h0);
    mcoreClass.set_mregs(32'h3eb, 32'h0);
    mcoreClass.set_mregs(32'h3ec, 32'h0);
    mcoreClass.set_mregs(32'h3ed, 32'h0);
    mcoreClass.set_mregs(32'h3ee, 32'h0);
    mcoreClass.set_mregs(32'h3ef, 32'h0);
    mcoreClass.set_mregs(32'h3f0, 32'h0);
    mcoreClass.set_mregs(32'h3f1, 32'h0);
    mcoreClass.set_mregs(32'h3f2, 32'h0);
    mcoreClass.set_mregs(32'h3f3, 32'h0);
    mcoreClass.set_mregs(32'h3f4, 32'h0);
    mcoreClass.set_mregs(32'h3f5, 32'h0);
    mcoreClass.set_mregs(32'h3f6, 32'h0);
    mcoreClass.set_mregs(32'h3f7, 32'h0);
    mcoreClass.set_mregs(32'h3f8, 32'h0);
    mcoreClass.set_mregs(32'h3f9, 32'h0);
    mcoreClass.set_mregs(32'h3fa, 32'h0);
    mcoreClass.set_mregs(32'h3fb, 32'h0);
    mcoreClass.set_mregs(32'h3fc, 32'h0);
    mcoreClass.set_mregs(32'h3fd, 32'h0);
    mcoreClass.set_mregs(32'h3fe, 32'h0);
    mcoreClass.set_mregs(32'h3ff, 32'h0);
    mcoreClass.set_mregs(32'h400, 32'h0);
    mcoreClass.set_mregs(32'h401, 32'h0);
    mcoreClass.set_mregs(32'h402, 32'h0);
    mcoreClass.set_mregs(32'h403, 32'h0);
    mcoreClass.set_mregs(32'h404, 32'h0);
    mcoreClass.set_mregs(32'h405, 32'h0);
    mcoreClass.set_mregs(32'h406, 32'h0);
    mcoreClass.set_mregs(32'h407, 32'h0);
    mcoreClass.set_mregs(32'h408, 32'h0);
    mcoreClass.set_mregs(32'h409, 32'h0);
    mcoreClass.set_mregs(32'h40a, 32'h0);
    mcoreClass.set_mregs(32'h40b, 32'h0);
    mcoreClass.set_mregs(32'h40c, 32'h0);
    mcoreClass.set_mregs(32'h40d, 32'h0);
    mcoreClass.set_mregs(32'h40e, 32'h0);
    mcoreClass.set_mregs(32'h40f, 32'h0);
    mcoreClass.set_mregs(32'h410, 32'h0);
    mcoreClass.set_mregs(32'h411, 32'h0);
    mcoreClass.set_mregs(32'h412, 32'h0);
    mcoreClass.set_mregs(32'h413, 32'h0);
    mcoreClass.set_mregs(32'h414, 32'h0);
    mcoreClass.set_mregs(32'h415, 32'h0);
    mcoreClass.set_mregs(32'h416, 32'h0);
    mcoreClass.set_mregs(32'h417, 32'h0);
    mcoreClass.set_mregs(32'h418, 32'h0);
    mcoreClass.set_mregs(32'h419, 32'h0);
    mcoreClass.set_mregs(32'h41a, 32'h0);
    mcoreClass.set_mregs(32'h41b, 32'h0);
    mcoreClass.set_mregs(32'h41c, 32'h0);
    mcoreClass.set_mregs(32'h41d, 32'h0);
    mcoreClass.set_mregs(32'h41e, 32'h0);
    mcoreClass.set_mregs(32'h41f, 32'h0);
    mcoreClass.set_mregs(32'h420, 32'h0);
    mcoreClass.set_mregs(32'h421, 32'h0);
    mcoreClass.set_mregs(32'h422, 32'h0);
    mcoreClass.set_mregs(32'h423, 32'h0);
    mcoreClass.set_mregs(32'h424, 32'h0);
    mcoreClass.set_mregs(32'h425, 32'h0);
    mcoreClass.set_mregs(32'h426, 32'h0);
    mcoreClass.set_mregs(32'h427, 32'h0);
    mcoreClass.set_mregs(32'h428, 32'h0);
    mcoreClass.set_mregs(32'h429, 32'h0);
    mcoreClass.set_mregs(32'h42a, 32'h0);
    mcoreClass.set_mregs(32'h42b, 32'h0);
    mcoreClass.set_mregs(32'h42c, 32'h0);
    mcoreClass.set_mregs(32'h42d, 32'h0);
    mcoreClass.set_mregs(32'h42e, 32'h0);
    mcoreClass.set_mregs(32'h42f, 32'h0);
    mcoreClass.set_mregs(32'h430, 32'h0);
    mcoreClass.set_mregs(32'h431, 32'h0);
    mcoreClass.set_mregs(32'h432, 32'h0);
    mcoreClass.set_mregs(32'h433, 32'h0);
    mcoreClass.set_mregs(32'h434, 32'h0);
    mcoreClass.set_mregs(32'h435, 32'h0);
    mcoreClass.set_mregs(32'h436, 32'h0);
    mcoreClass.set_mregs(32'h437, 32'h0);
    mcoreClass.set_mregs(32'h438, 32'h0);
    mcoreClass.set_mregs(32'h439, 32'h0);
    mcoreClass.set_mregs(32'h43a, 32'h0);
    mcoreClass.set_mregs(32'h43b, 32'h0);
    mcoreClass.set_mregs(32'h43c, 32'h0);
    mcoreClass.set_mregs(32'h43d, 32'h0);
    mcoreClass.set_mregs(32'h43e, 32'h0);
    mcoreClass.set_mregs(32'h43f, 32'h0);
    mcoreClass.set_mregs(32'h440, 32'h0);
    mcoreClass.set_mregs(32'h441, 32'h0);
    mcoreClass.set_mregs(32'h442, 32'h0);
    mcoreClass.set_mregs(32'h443, 32'h0);
    mcoreClass.set_mregs(32'h444, 32'h0);
    mcoreClass.set_mregs(32'h445, 32'h0);
    mcoreClass.set_mregs(32'h446, 32'h0);
    mcoreClass.set_mregs(32'h447, 32'h0);
    mcoreClass.set_mregs(32'h448, 32'h0);
    mcoreClass.set_mregs(32'h449, 32'h0);
    mcoreClass.set_mregs(32'h44a, 32'h0);
    mcoreClass.set_mregs(32'h44b, 32'h0);
    mcoreClass.set_mregs(32'h44c, 32'h0);
    mcoreClass.set_mregs(32'h44d, 32'h0);
    mcoreClass.set_mregs(32'h44e, 32'h0);
    mcoreClass.set_mregs(32'h44f, 32'h0);
    mcoreClass.set_mregs(32'h450, 32'h0);
    mcoreClass.set_mregs(32'h451, 32'h0);
    mcoreClass.set_mregs(32'h452, 32'h0);
    mcoreClass.set_mregs(32'h453, 32'h0);
    mcoreClass.set_mregs(32'h454, 32'h0);
    mcoreClass.set_mregs(32'h455, 32'h0);
    mcoreClass.set_mregs(32'h456, 32'h0);
    mcoreClass.set_mregs(32'h457, 32'h0);
    mcoreClass.set_mregs(32'h458, 32'h0);
    mcoreClass.set_mregs(32'h459, 32'h0);
    mcoreClass.set_mregs(32'h45a, 32'h0);
    mcoreClass.set_mregs(32'h45b, 32'h0);
    mcoreClass.set_mregs(32'h45c, 32'h0);
    mcoreClass.set_mregs(32'h45d, 32'h0);
    mcoreClass.set_mregs(32'h45e, 32'h0);
    mcoreClass.set_mregs(32'h45f, 32'h0);
    mcoreClass.set_mregs(32'h460, 32'h0);
    mcoreClass.set_mregs(32'h461, 32'h0);
    mcoreClass.set_mregs(32'h462, 32'h0);
    mcoreClass.set_mregs(32'h463, 32'h0);
    mcoreClass.set_mregs(32'h464, 32'h0);
    mcoreClass.set_mregs(32'h465, 32'h0);
    mcoreClass.set_mregs(32'h466, 32'h0);
    mcoreClass.set_mregs(32'h467, 32'h0);
    mcoreClass.set_mregs(32'h468, 32'h0);
    mcoreClass.set_mregs(32'h469, 32'h0);
    mcoreClass.set_mregs(32'h46a, 32'h0);
    mcoreClass.set_mregs(32'h46b, 32'h0);
    mcoreClass.set_mregs(32'h46c, 32'h0);
    mcoreClass.set_mregs(32'h46d, 32'h0);
    mcoreClass.set_mregs(32'h46e, 32'h0);
    mcoreClass.set_mregs(32'h46f, 32'h0);
    mcoreClass.set_mregs(32'h470, 32'h0);
    mcoreClass.set_mregs(32'h471, 32'h0);
    mcoreClass.set_mregs(32'h472, 32'h0);
    mcoreClass.set_mregs(32'h473, 32'h0);
    mcoreClass.set_mregs(32'h474, 32'h0);
    mcoreClass.set_mregs(32'h475, 32'h0);
    mcoreClass.set_mregs(32'h476, 32'h0);
    mcoreClass.set_mregs(32'h477, 32'h0);
    mcoreClass.set_mregs(32'h478, 32'h0);
    mcoreClass.set_mregs(32'h479, 32'h0);
    mcoreClass.set_mregs(32'h47a, 32'h0);
    mcoreClass.set_mregs(32'h47b, 32'h0);
    mcoreClass.set_mregs(32'h47c, 32'h0);
    mcoreClass.set_mregs(32'h47d, 32'h0);
    mcoreClass.set_mregs(32'h47e, 32'h0);
    mcoreClass.set_mregs(32'h47f, 32'h0);
    mcoreClass.set_mregs(32'h480, 32'h0);
    mcoreClass.set_mregs(32'h481, 32'h0);
    mcoreClass.set_mregs(32'h482, 32'h0);
    mcoreClass.set_mregs(32'h483, 32'h0);
    mcoreClass.set_mregs(32'h484, 32'h0);
    mcoreClass.set_mregs(32'h485, 32'h0);
    mcoreClass.set_mregs(32'h486, 32'h0);
    mcoreClass.set_mregs(32'h487, 32'h0);
    mcoreClass.set_mregs(32'h488, 32'h0);
    mcoreClass.set_mregs(32'h489, 32'h0);
    mcoreClass.set_mregs(32'h48a, 32'h0);
    mcoreClass.set_mregs(32'h48b, 32'h0);
    mcoreClass.set_mregs(32'h48c, 32'h0);
    mcoreClass.set_mregs(32'h48d, 32'h0);
    mcoreClass.set_mregs(32'h48e, 32'h0);
    mcoreClass.set_mregs(32'h48f, 32'h0);
    mcoreClass.set_mregs(32'h490, 32'h0);
    mcoreClass.set_mregs(32'h491, 32'h0);
    mcoreClass.set_mregs(32'h492, 32'h0);
    mcoreClass.set_mregs(32'h493, 32'h0);
    mcoreClass.set_mregs(32'h494, 32'h0);
    mcoreClass.set_mregs(32'h495, 32'h0);
    mcoreClass.set_mregs(32'h496, 32'h0);
    mcoreClass.set_mregs(32'h497, 32'h0);
    mcoreClass.set_mregs(32'h498, 32'h0);
    mcoreClass.set_mregs(32'h499, 32'h0);
    mcoreClass.set_mregs(32'h49a, 32'h0);
    mcoreClass.set_mregs(32'h49b, 32'h0);
    mcoreClass.set_mregs(32'h49c, 32'h0);
    mcoreClass.set_mregs(32'h49d, 32'h0);
    mcoreClass.set_mregs(32'h49e, 32'h0);
    mcoreClass.set_mregs(32'h49f, 32'h0);
    mcoreClass.set_mregs(32'h4a0, 32'h0);
    mcoreClass.set_mregs(32'h4a1, 32'h0);
    mcoreClass.set_mregs(32'h4a2, 32'h0);
    mcoreClass.set_mregs(32'h4a3, 32'h0);
    mcoreClass.set_mregs(32'h4a4, 32'h0);
    mcoreClass.set_mregs(32'h4a5, 32'h0);
    mcoreClass.set_mregs(32'h4a6, 32'h0);
    mcoreClass.set_mregs(32'h4a7, 32'h0);
    mcoreClass.set_mregs(32'h4a8, 32'h0);
    mcoreClass.set_mregs(32'h4a9, 32'h0);
    mcoreClass.set_mregs(32'h4aa, 32'h0);
    mcoreClass.set_mregs(32'h4ab, 32'h0);
    mcoreClass.set_mregs(32'h4ac, 32'h0);
    mcoreClass.set_mregs(32'h4ad, 32'h0);
    mcoreClass.set_mregs(32'h4ae, 32'h0);
    mcoreClass.set_mregs(32'h4af, 32'h0);
    mcoreClass.set_mregs(32'h4b0, 32'h0);
    mcoreClass.set_mregs(32'h4b1, 32'h0);
    mcoreClass.set_mregs(32'h4b2, 32'h0);
    mcoreClass.set_mregs(32'h4b3, 32'h0);
    mcoreClass.set_mregs(32'h4b4, 32'h0);
    mcoreClass.set_mregs(32'h4b5, 32'h0);
    mcoreClass.set_mregs(32'h4b6, 32'h0);
    mcoreClass.set_mregs(32'h4b7, 32'h0);
    mcoreClass.set_mregs(32'h4b8, 32'h0);
    mcoreClass.set_mregs(32'h4b9, 32'h0);
    mcoreClass.set_mregs(32'h4ba, 32'h0);
    mcoreClass.set_mregs(32'h4bb, 32'h0);
    mcoreClass.set_mregs(32'h4bc, 32'h0);
    mcoreClass.set_mregs(32'h4bd, 32'h0);
    mcoreClass.set_mregs(32'h4be, 32'h0);
    mcoreClass.set_mregs(32'h4bf, 32'h0);
    mcoreClass.set_mregs(32'h4c0, 32'h0);
    mcoreClass.set_mregs(32'h4c1, 32'h0);
    mcoreClass.set_mregs(32'h4c2, 32'h0);
    mcoreClass.set_mregs(32'h4c3, 32'h0);
    mcoreClass.set_mregs(32'h4c4, 32'h0);
    mcoreClass.set_mregs(32'h4c5, 32'h0);
    mcoreClass.set_mregs(32'h4c6, 32'h0);
    mcoreClass.set_mregs(32'h4c7, 32'h0);
    mcoreClass.set_mregs(32'h4c8, 32'h0);
    mcoreClass.set_mregs(32'h4c9, 32'h0);
    mcoreClass.set_mregs(32'h4ca, 32'h0);
    mcoreClass.set_mregs(32'h4cb, 32'h0);
    mcoreClass.set_mregs(32'h4cc, 32'h0);
    mcoreClass.set_mregs(32'h4cd, 32'h0);
    mcoreClass.set_mregs(32'h4ce, 32'h0);
    mcoreClass.set_mregs(32'h4cf, 32'h0);
    mcoreClass.set_mregs(32'h4d0, 32'h0);
    mcoreClass.set_mregs(32'h4d1, 32'h0);
    mcoreClass.set_mregs(32'h4d2, 32'h0);
    mcoreClass.set_mregs(32'h4d3, 32'h0);
    mcoreClass.set_mregs(32'h4d4, 32'h0);
    mcoreClass.set_mregs(32'h4d5, 32'h0);
    mcoreClass.set_mregs(32'h4d6, 32'h0);
    mcoreClass.set_mregs(32'h4d7, 32'h0);
    mcoreClass.set_mregs(32'h4d8, 32'h0);
    mcoreClass.set_mregs(32'h4d9, 32'h0);
    mcoreClass.set_mregs(32'h4da, 32'h0);
    mcoreClass.set_mregs(32'h4db, 32'h0);
    mcoreClass.set_mregs(32'h4dc, 32'h0);
    mcoreClass.set_mregs(32'h4dd, 32'h0);
    mcoreClass.set_mregs(32'h4de, 32'h0);
    mcoreClass.set_mregs(32'h4df, 32'h0);
    mcoreClass.set_mregs(32'h4e0, 32'h0);
    mcoreClass.set_mregs(32'h4e1, 32'h0);
    mcoreClass.set_mregs(32'h4e2, 32'h0);
    mcoreClass.set_mregs(32'h4e3, 32'h0);
    mcoreClass.set_mregs(32'h4e4, 32'h0);
    mcoreClass.set_mregs(32'h4e5, 32'h0);
    mcoreClass.set_mregs(32'h4e6, 32'h0);
    mcoreClass.set_mregs(32'h4e7, 32'h0);
    mcoreClass.set_mregs(32'h4e8, 32'h0);
    mcoreClass.set_mregs(32'h4e9, 32'h0);
    mcoreClass.set_mregs(32'h4ea, 32'h0);
    mcoreClass.set_mregs(32'h4eb, 32'h0);
    mcoreClass.set_mregs(32'h4ec, 32'h0);
    mcoreClass.set_mregs(32'h4ed, 32'h0);
    mcoreClass.set_mregs(32'h4ee, 32'h0);
    mcoreClass.set_mregs(32'h4ef, 32'h0);
    mcoreClass.set_mregs(32'h4f0, 32'h0);
    mcoreClass.set_mregs(32'h4f1, 32'h0);
    mcoreClass.set_mregs(32'h4f2, 32'h0);
    mcoreClass.set_mregs(32'h4f3, 32'h0);
    mcoreClass.set_mregs(32'h4f4, 32'h0);
    mcoreClass.set_mregs(32'h4f5, 32'h0);
    mcoreClass.set_mregs(32'h4f6, 32'h0);
    mcoreClass.set_mregs(32'h4f7, 32'h0);
    mcoreClass.set_mregs(32'h4f8, 32'h0);
    mcoreClass.set_mregs(32'h4f9, 32'h0);
    mcoreClass.set_mregs(32'h4fa, 32'h0);
    mcoreClass.set_mregs(32'h4fb, 32'h0);
    mcoreClass.set_mregs(32'h4fc, 32'h0);
    mcoreClass.set_mregs(32'h4fd, 32'h0);
    mcoreClass.set_mregs(32'h4fe, 32'h0);
    mcoreClass.set_mregs(32'h4ff, 32'h0);
    mcoreClass.set_mregs(32'h500, 32'h0);
    mcoreClass.set_mregs(32'h501, 32'h0);
    mcoreClass.set_mregs(32'h502, 32'h0);
    mcoreClass.set_mregs(32'h503, 32'h0);
    mcoreClass.set_mregs(32'h504, 32'h0);
    mcoreClass.set_mregs(32'h505, 32'h0);
    mcoreClass.set_mregs(32'h506, 32'h0);
    mcoreClass.set_mregs(32'h507, 32'h0);
    mcoreClass.set_mregs(32'h508, 32'h0);
    mcoreClass.set_mregs(32'h509, 32'h0);
    mcoreClass.set_mregs(32'h50a, 32'h0);
    mcoreClass.set_mregs(32'h50b, 32'h0);
    mcoreClass.set_mregs(32'h50c, 32'h0);
    mcoreClass.set_mregs(32'h50d, 32'h0);
    mcoreClass.set_mregs(32'h50e, 32'h0);
    mcoreClass.set_mregs(32'h50f, 32'h0);
    mcoreClass.set_mregs(32'h510, 32'h0);
    mcoreClass.set_mregs(32'h511, 32'h0);
    mcoreClass.set_mregs(32'h512, 32'h0);
    mcoreClass.set_mregs(32'h513, 32'h0);
    mcoreClass.set_mregs(32'h514, 32'h0);
    mcoreClass.set_mregs(32'h515, 32'h0);
    mcoreClass.set_mregs(32'h516, 32'h0);
    mcoreClass.set_mregs(32'h517, 32'h0);
    mcoreClass.set_mregs(32'h518, 32'h0);
    mcoreClass.set_mregs(32'h519, 32'h0);
    mcoreClass.set_mregs(32'h51a, 32'h0);
    mcoreClass.set_mregs(32'h51b, 32'h0);
    mcoreClass.set_mregs(32'h51c, 32'h0);
    mcoreClass.set_mregs(32'h51d, 32'h0);
    mcoreClass.set_mregs(32'h51e, 32'h0);
    mcoreClass.set_mregs(32'h51f, 32'h0);
    mcoreClass.set_mregs(32'h520, 32'h0);
    mcoreClass.set_mregs(32'h521, 32'h0);
    mcoreClass.set_mregs(32'h522, 32'h0);
    mcoreClass.set_mregs(32'h523, 32'h0);
    mcoreClass.set_mregs(32'h524, 32'h0);
    mcoreClass.set_mregs(32'h525, 32'h0);
    mcoreClass.set_mregs(32'h526, 32'h0);
    mcoreClass.set_mregs(32'h527, 32'h0);
    mcoreClass.set_mregs(32'h528, 32'h0);
    mcoreClass.set_mregs(32'h529, 32'h0);
    mcoreClass.set_mregs(32'h52a, 32'h0);
    mcoreClass.set_mregs(32'h52b, 32'h0);
    mcoreClass.set_mregs(32'h52c, 32'h0);
    mcoreClass.set_mregs(32'h52d, 32'h0);
    mcoreClass.set_mregs(32'h52e, 32'h0);
    mcoreClass.set_mregs(32'h52f, 32'h0);
    mcoreClass.set_mregs(32'h530, 32'h0);
    mcoreClass.set_mregs(32'h531, 32'h0);
    mcoreClass.set_mregs(32'h532, 32'h0);
    mcoreClass.set_mregs(32'h533, 32'h0);
    mcoreClass.set_mregs(32'h534, 32'h0);
    mcoreClass.set_mregs(32'h535, 32'h0);
    mcoreClass.set_mregs(32'h536, 32'h0);
    mcoreClass.set_mregs(32'h537, 32'h0);
    mcoreClass.set_mregs(32'h538, 32'h0);
    mcoreClass.set_mregs(32'h539, 32'h0);
    mcoreClass.set_mregs(32'h53a, 32'h0);
    mcoreClass.set_mregs(32'h53b, 32'h0);
    mcoreClass.set_mregs(32'h53c, 32'h0);
    mcoreClass.set_mregs(32'h53d, 32'h0);
    mcoreClass.set_mregs(32'h53e, 32'h0);
    mcoreClass.set_mregs(32'h53f, 32'h0);
    mcoreClass.set_mregs(32'h540, 32'h251b7c);
    mcoreClass.set_mregs(32'h541, 32'h0);
    mcoreClass.set_mregs(32'h542, 32'h0);
    mcoreClass.set_mregs(32'h543, 32'h0);
    mcoreClass.set_mregs(32'h544, 32'hfffffffc);
    mcoreClass.set_mregs(32'h545, 32'h0);
    mcoreClass.set_mregs(32'h546, 32'h0);
    mcoreClass.set_mregs(32'h547, 32'h0);
    mcoreClass.set_mregs(32'h548, 32'h0);
    mcoreClass.set_mregs(32'h549, 32'h0);
    mcoreClass.set_mregs(32'h54a, 32'h0);
    mcoreClass.set_mregs(32'h54b, 32'h0);
    mcoreClass.set_mregs(32'h54c, 32'h0);
    mcoreClass.set_mregs(32'h54d, 32'h0);
    mcoreClass.set_mregs(32'h54e, 32'h0);
    mcoreClass.set_mregs(32'h54f, 32'h0);
    mcoreClass.set_mregs(32'h550, 32'h0);
    mcoreClass.set_mregs(32'h551, 32'h0);
    mcoreClass.set_mregs(32'h552, 32'h0);
    mcoreClass.set_mregs(32'h553, 32'h0);
    mcoreClass.set_mregs(32'h554, 32'h0);
    mcoreClass.set_mregs(32'h555, 32'h0);
    mcoreClass.set_mregs(32'h556, 32'h0);
    mcoreClass.set_mregs(32'h557, 32'h0);
    mcoreClass.set_mregs(32'h558, 32'h0);
    mcoreClass.set_mregs(32'h559, 32'h0);
    mcoreClass.set_mregs(32'h55a, 32'h0);
    mcoreClass.set_mregs(32'h55b, 32'h0);
    mcoreClass.set_mregs(32'h55c, 32'h0);
    mcoreClass.set_mregs(32'h55d, 32'h0);
    mcoreClass.set_mregs(32'h55e, 32'h0);
    mcoreClass.set_mregs(32'h55f, 32'h0);
    mcoreClass.set_mregs(32'h560, 32'h0);
    mcoreClass.set_mregs(32'h561, 32'h0);
    mcoreClass.set_mregs(32'h562, 32'h0);
    mcoreClass.set_mregs(32'h563, 32'h0);
    mcoreClass.set_mregs(32'h564, 32'h0);
    mcoreClass.set_mregs(32'h565, 32'h0);
    mcoreClass.set_mregs(32'h566, 32'h0);
    mcoreClass.set_mregs(32'h567, 32'h0);
    mcoreClass.set_mregs(32'h568, 32'h0);
    mcoreClass.set_mregs(32'h569, 32'h0);
    mcoreClass.set_mregs(32'h56a, 32'h0);
    mcoreClass.set_mregs(32'h56b, 32'h0);
    mcoreClass.set_mregs(32'h56c, 32'h0);
    mcoreClass.set_mregs(32'h56d, 32'h0);
    mcoreClass.set_mregs(32'h56e, 32'h0);
    mcoreClass.set_mregs(32'h56f, 32'h0);
    mcoreClass.set_mregs(32'h570, 32'h1fcc04);
    mcoreClass.set_mregs(32'h571, 32'h0);
    mcoreClass.set_mregs(32'h572, 32'h0);
    mcoreClass.set_mregs(32'h573, 32'h0);
    mcoreClass.set_mregs(32'h574, 32'hfffffffc);
    mcoreClass.set_mregs(32'h575, 32'h0);
    mcoreClass.set_mregs(32'h576, 32'h0);
    mcoreClass.set_mregs(32'h577, 32'h0);
    mcoreClass.set_mregs(32'h578, 32'h1fcb34);
    mcoreClass.set_mregs(32'h579, 32'h0);
    mcoreClass.set_mregs(32'h57a, 32'h0);
    mcoreClass.set_mregs(32'h57b, 32'h0);
    mcoreClass.set_mregs(32'h57c, 32'h0);
    mcoreClass.set_mregs(32'h57d, 32'h0);
    mcoreClass.set_mregs(32'h57e, 32'h0);
    mcoreClass.set_mregs(32'h57f, 32'h0);
    mcoreClass.set_mregs(32'h580, 32'h0);
    mcoreClass.set_mregs(32'h581, 32'h0);
    mcoreClass.set_mregs(32'h582, 32'h0);
    mcoreClass.set_mregs(32'h583, 32'h0);
    mcoreClass.set_mregs(32'h584, 32'h0);
    mcoreClass.set_mregs(32'h585, 32'h0);
    mcoreClass.set_mregs(32'h586, 32'h0);
    mcoreClass.set_mregs(32'h587, 32'h0);
    mcoreClass.set_mregs(32'h588, 32'h0);
    mcoreClass.set_mregs(32'h589, 32'h0);
    mcoreClass.set_mregs(32'h58a, 32'h0);
    mcoreClass.set_mregs(32'h58b, 32'h0);
    mcoreClass.set_mregs(32'h58c, 32'h0);
    mcoreClass.set_mregs(32'h58d, 32'h0);
    mcoreClass.set_mregs(32'h58e, 32'h0);
    mcoreClass.set_mregs(32'h58f, 32'h0);
    mcoreClass.set_mregs(32'h590, 32'h0);
    mcoreClass.set_mregs(32'h591, 32'h0);
    mcoreClass.set_mregs(32'h592, 32'h0);
    mcoreClass.set_mregs(32'h593, 32'h0);
    mcoreClass.set_mregs(32'h594, 32'h0);
    mcoreClass.set_mregs(32'h595, 32'h0);
    mcoreClass.set_mregs(32'h596, 32'h0);
    mcoreClass.set_mregs(32'h597, 32'h0);
    mcoreClass.set_mregs(32'h598, 32'h0);
    mcoreClass.set_mregs(32'h599, 32'h0);
    mcoreClass.set_mregs(32'h59a, 32'h0);
    mcoreClass.set_mregs(32'h59b, 32'h0);
    mcoreClass.set_mregs(32'h59c, 32'h0);
    mcoreClass.set_mregs(32'h59d, 32'h0);
    mcoreClass.set_mregs(32'h59e, 32'h0);
    mcoreClass.set_mregs(32'h59f, 32'h0);
    mcoreClass.set_mregs(32'h5a0, 32'h1006d0);
    mcoreClass.set_mregs(32'h5a1, 32'h0);
    mcoreClass.set_mregs(32'h5a2, 32'h0);
    mcoreClass.set_mregs(32'h5a3, 32'h0);
    mcoreClass.set_mregs(32'h5a4, 32'h1006d0);
    mcoreClass.set_mregs(32'h5a5, 32'h0);
    mcoreClass.set_mregs(32'h5a6, 32'h0);
    mcoreClass.set_mregs(32'h5a7, 32'h0);
    mcoreClass.set_mregs(32'h5a8, 32'h28db50);
    mcoreClass.set_mregs(32'h5a9, 32'h0);
    mcoreClass.set_mregs(32'h5aa, 32'h0);
    mcoreClass.set_mregs(32'h5ab, 32'h0);
    mcoreClass.set_mregs(32'h5ac, 32'h283b08);
    mcoreClass.set_mregs(32'h5ad, 32'h0);
    mcoreClass.set_mregs(32'h5ae, 32'h0);
    mcoreClass.set_mregs(32'h5af, 32'h0);
    mcoreClass.set_mregs(32'h5b0, 32'h0);
    mcoreClass.set_mregs(32'h5b1, 32'h0);
    mcoreClass.set_mregs(32'h5b2, 32'h0);
    mcoreClass.set_mregs(32'h5b3, 32'h0);
    mcoreClass.set_mregs(32'h5b4, 32'h0);
    mcoreClass.set_mregs(32'h5b5, 32'h0);
    mcoreClass.set_mregs(32'h5b6, 32'h0);
    mcoreClass.set_mregs(32'h5b7, 32'h0);
    mcoreClass.set_mregs(32'h5b8, 32'h0);
    mcoreClass.set_mregs(32'h5b9, 32'h0);
    mcoreClass.set_mregs(32'h5ba, 32'h0);
    mcoreClass.set_mregs(32'h5bb, 32'h0);
    mcoreClass.set_mregs(32'h5bc, 32'h0);
    mcoreClass.set_mregs(32'h5bd, 32'h0);
    mcoreClass.set_mregs(32'h5be, 32'h0);
    mcoreClass.set_mregs(32'h5bf, 32'h0);
    mcoreClass.set_mregs(32'h5c0, 32'h0);
    mcoreClass.set_mregs(32'h5c1, 32'h0);
    mcoreClass.set_mregs(32'h5c2, 32'h0);
    mcoreClass.set_mregs(32'h5c3, 32'h0);
    mcoreClass.set_mregs(32'h5c4, 32'h0);
    mcoreClass.set_mregs(32'h5c5, 32'h0);
    mcoreClass.set_mregs(32'h5c6, 32'h0);
    mcoreClass.set_mregs(32'h5c7, 32'h0);
    mcoreClass.set_mregs(32'h5c8, 32'h0);
    mcoreClass.set_mregs(32'h5c9, 32'h0);
    mcoreClass.set_mregs(32'h5ca, 32'h0);
    mcoreClass.set_mregs(32'h5cb, 32'h0);
    mcoreClass.set_mregs(32'h5cc, 32'h0);
    mcoreClass.set_mregs(32'h5cd, 32'h0);
    mcoreClass.set_mregs(32'h5ce, 32'h0);
    mcoreClass.set_mregs(32'h5cf, 32'h0);
    mcoreClass.set_mregs(32'h5d0, 32'h0);
    mcoreClass.set_mregs(32'h5d1, 32'h0);
    mcoreClass.set_mregs(32'h5d2, 32'h0);
    mcoreClass.set_mregs(32'h5d3, 32'h0);
    mcoreClass.set_mregs(32'h5d4, 32'h0);
    mcoreClass.set_mregs(32'h5d5, 32'h0);
    mcoreClass.set_mregs(32'h5d6, 32'h0);
    mcoreClass.set_mregs(32'h5d7, 32'h0);
    mcoreClass.set_mregs(32'h5d8, 32'h0);
    mcoreClass.set_mregs(32'h5d9, 32'h0);
    mcoreClass.set_mregs(32'h5da, 32'h0);
    mcoreClass.set_mregs(32'h5db, 32'h0);
    mcoreClass.set_mregs(32'h5dc, 32'h0);
    mcoreClass.set_mregs(32'h5dd, 32'h0);
    mcoreClass.set_mregs(32'h5de, 32'h0);
    mcoreClass.set_mregs(32'h5df, 32'h0);
    mcoreClass.set_mregs(32'h5e0, 32'h0);
    mcoreClass.set_mregs(32'h5e1, 32'h0);
    mcoreClass.set_mregs(32'h5e2, 32'h0);
    mcoreClass.set_mregs(32'h5e3, 32'h0);
    mcoreClass.set_mregs(32'h5e4, 32'h0);
    mcoreClass.set_mregs(32'h5e5, 32'h0);
    mcoreClass.set_mregs(32'h5e6, 32'h0);
    mcoreClass.set_mregs(32'h5e7, 32'h0);
    mcoreClass.set_mregs(32'h5e8, 32'h0);
    mcoreClass.set_mregs(32'h5e9, 32'h0);
    mcoreClass.set_mregs(32'h5ea, 32'h0);
    mcoreClass.set_mregs(32'h5eb, 32'h0);
    mcoreClass.set_mregs(32'h5ec, 32'h0);
    mcoreClass.set_mregs(32'h5ed, 32'h0);
    mcoreClass.set_mregs(32'h5ee, 32'h0);
    mcoreClass.set_mregs(32'h5ef, 32'h0);
    mcoreClass.set_mregs(32'h5f0, 32'h0);
    mcoreClass.set_mregs(32'h5f1, 32'h0);
    mcoreClass.set_mregs(32'h5f2, 32'h0);
    mcoreClass.set_mregs(32'h5f3, 32'h0);
    mcoreClass.set_mregs(32'h5f4, 32'h0);
    mcoreClass.set_mregs(32'h5f5, 32'h0);
    mcoreClass.set_mregs(32'h5f6, 32'h0);
    mcoreClass.set_mregs(32'h5f7, 32'h0);
    mcoreClass.set_mregs(32'h5f8, 32'h0);
    mcoreClass.set_mregs(32'h5f9, 32'h0);
    mcoreClass.set_mregs(32'h5fa, 32'h0);
    mcoreClass.set_mregs(32'h5fb, 32'h0);
    mcoreClass.set_mregs(32'h5fc, 32'h0);
    mcoreClass.set_mregs(32'h5fd, 32'h0);
    mcoreClass.set_mregs(32'h5fe, 32'h0);
    mcoreClass.set_mregs(32'h5ff, 32'h0);
    mcoreClass.set_mregs(32'h600, 32'h0);
    mcoreClass.set_mregs(32'h601, 32'h0);
    mcoreClass.set_mregs(32'h602, 32'h0);
    mcoreClass.set_mregs(32'h603, 32'h0);
    mcoreClass.set_mregs(32'h604, 32'h0);
    mcoreClass.set_mregs(32'h605, 32'h0);
    mcoreClass.set_mregs(32'h606, 32'h0);
    mcoreClass.set_mregs(32'h607, 32'h0);
    mcoreClass.set_mregs(32'h608, 32'h0);
    mcoreClass.set_mregs(32'h609, 32'h0);
    mcoreClass.set_mregs(32'h60a, 32'h0);
    mcoreClass.set_mregs(32'h60b, 32'h0);
    mcoreClass.set_mregs(32'h60c, 32'h0);
    mcoreClass.set_mregs(32'h60d, 32'h0);
    mcoreClass.set_mregs(32'h60e, 32'h0);
    mcoreClass.set_mregs(32'h60f, 32'h0);
    mcoreClass.set_mregs(32'h610, 32'h0);
    mcoreClass.set_mregs(32'h611, 32'h0);
    mcoreClass.set_mregs(32'h612, 32'h0);
    mcoreClass.set_mregs(32'h613, 32'h0);
    mcoreClass.set_mregs(32'h614, 32'h0);
    mcoreClass.set_mregs(32'h615, 32'h0);
    mcoreClass.set_mregs(32'h616, 32'h0);
    mcoreClass.set_mregs(32'h617, 32'h0);
    mcoreClass.set_mregs(32'h618, 32'h0);
    mcoreClass.set_mregs(32'h619, 32'h0);
    mcoreClass.set_mregs(32'h61a, 32'h0);
    mcoreClass.set_mregs(32'h61b, 32'h0);
    mcoreClass.set_mregs(32'h61c, 32'h0);
    mcoreClass.set_mregs(32'h61d, 32'h0);
    mcoreClass.set_mregs(32'h61e, 32'h0);
    mcoreClass.set_mregs(32'h61f, 32'h0);
    mcoreClass.set_mregs(32'h620, 32'h0);
    mcoreClass.set_mregs(32'h621, 32'h0);
    mcoreClass.set_mregs(32'h622, 32'h0);
    mcoreClass.set_mregs(32'h623, 32'h0);
    mcoreClass.set_mregs(32'h624, 32'h0);
    mcoreClass.set_mregs(32'h625, 32'h0);
    mcoreClass.set_mregs(32'h626, 32'h0);
    mcoreClass.set_mregs(32'h627, 32'h0);
    mcoreClass.set_mregs(32'h628, 32'h0);
    mcoreClass.set_mregs(32'h629, 32'h0);
    mcoreClass.set_mregs(32'h62a, 32'h0);
    mcoreClass.set_mregs(32'h62b, 32'h0);
    mcoreClass.set_mregs(32'h62c, 32'h0);
    mcoreClass.set_mregs(32'h62d, 32'h0);
    mcoreClass.set_mregs(32'h62e, 32'h0);
    mcoreClass.set_mregs(32'h62f, 32'h0);
    mcoreClass.set_mregs(32'h630, 32'h0);
    mcoreClass.set_mregs(32'h631, 32'h0);
    mcoreClass.set_mregs(32'h632, 32'h0);
    mcoreClass.set_mregs(32'h633, 32'h0);
    mcoreClass.set_mregs(32'h634, 32'h0);
    mcoreClass.set_mregs(32'h635, 32'h0);
    mcoreClass.set_mregs(32'h636, 32'h0);
    mcoreClass.set_mregs(32'h637, 32'h0);
    mcoreClass.set_mregs(32'h638, 32'h0);
    mcoreClass.set_mregs(32'h639, 32'h0);
    mcoreClass.set_mregs(32'h63a, 32'h0);
    mcoreClass.set_mregs(32'h63b, 32'h0);
    mcoreClass.set_mregs(32'h63c, 32'h0);
    mcoreClass.set_mregs(32'h63d, 32'h0);
    mcoreClass.set_mregs(32'h63e, 32'h0);
    mcoreClass.set_mregs(32'h63f, 32'h0);
    mcoreClass.set_mregs(32'h640, 32'h0);
    mcoreClass.set_mregs(32'h641, 32'h0);
    mcoreClass.set_mregs(32'h642, 32'h0);
    mcoreClass.set_mregs(32'h643, 32'h0);
    mcoreClass.set_mregs(32'h644, 32'h0);
    mcoreClass.set_mregs(32'h645, 32'h0);
    mcoreClass.set_mregs(32'h646, 32'h0);
    mcoreClass.set_mregs(32'h647, 32'h0);
    mcoreClass.set_mregs(32'h648, 32'h0);
    mcoreClass.set_mregs(32'h649, 32'h0);
    mcoreClass.set_mregs(32'h64a, 32'h0);
    mcoreClass.set_mregs(32'h64b, 32'h0);
    mcoreClass.set_mregs(32'h64c, 32'h0);
    mcoreClass.set_mregs(32'h64d, 32'h0);
    mcoreClass.set_mregs(32'h64e, 32'h0);
    mcoreClass.set_mregs(32'h64f, 32'h0);
    mcoreClass.set_mregs(32'h650, 32'h0);
    mcoreClass.set_mregs(32'h651, 32'h0);
    mcoreClass.set_mregs(32'h652, 32'h0);
    mcoreClass.set_mregs(32'h653, 32'h0);
    mcoreClass.set_mregs(32'h654, 32'h0);
    mcoreClass.set_mregs(32'h655, 32'h0);
    mcoreClass.set_mregs(32'h656, 32'h0);
    mcoreClass.set_mregs(32'h657, 32'h0);
    mcoreClass.set_mregs(32'h658, 32'h0);
    mcoreClass.set_mregs(32'h659, 32'h0);
    mcoreClass.set_mregs(32'h65a, 32'h0);
    mcoreClass.set_mregs(32'h65b, 32'h0);
    mcoreClass.set_mregs(32'h65c, 32'h0);
    mcoreClass.set_mregs(32'h65d, 32'h0);
    mcoreClass.set_mregs(32'h65e, 32'h0);
    mcoreClass.set_mregs(32'h65f, 32'h0);
    mcoreClass.set_mregs(32'h660, 32'h0);
    mcoreClass.set_mregs(32'h661, 32'h0);
    mcoreClass.set_mregs(32'h662, 32'h0);
    mcoreClass.set_mregs(32'h663, 32'h0);
    mcoreClass.set_mregs(32'h664, 32'h0);
    mcoreClass.set_mregs(32'h665, 32'h0);
    mcoreClass.set_mregs(32'h666, 32'h0);
    mcoreClass.set_mregs(32'h667, 32'h0);
    mcoreClass.set_mregs(32'h668, 32'h0);
    mcoreClass.set_mregs(32'h669, 32'h0);
    mcoreClass.set_mregs(32'h66a, 32'h0);
    mcoreClass.set_mregs(32'h66b, 32'h0);
    mcoreClass.set_mregs(32'h66c, 32'h0);
    mcoreClass.set_mregs(32'h66d, 32'h0);
    mcoreClass.set_mregs(32'h66e, 32'h0);
    mcoreClass.set_mregs(32'h66f, 32'h0);
    mcoreClass.set_mregs(32'h670, 32'h0);
    mcoreClass.set_mregs(32'h671, 32'h0);
    mcoreClass.set_mregs(32'h672, 32'h0);
    mcoreClass.set_mregs(32'h673, 32'h0);
    mcoreClass.set_mregs(32'h674, 32'h0);
    mcoreClass.set_mregs(32'h675, 32'h0);
    mcoreClass.set_mregs(32'h676, 32'h0);
    mcoreClass.set_mregs(32'h677, 32'h0);
    mcoreClass.set_mregs(32'h678, 32'h0);
    mcoreClass.set_mregs(32'h679, 32'h0);
    mcoreClass.set_mregs(32'h67a, 32'h0);
    mcoreClass.set_mregs(32'h67b, 32'h0);
    mcoreClass.set_mregs(32'h67c, 32'h0);
    mcoreClass.set_mregs(32'h67d, 32'h0);
    mcoreClass.set_mregs(32'h67e, 32'h0);
    mcoreClass.set_mregs(32'h67f, 32'h0);
    mcoreClass.set_mregs(32'h680, 32'h0);
    mcoreClass.set_mregs(32'h681, 32'h0);
    mcoreClass.set_mregs(32'h682, 32'h0);
    mcoreClass.set_mregs(32'h683, 32'h0);
    mcoreClass.set_mregs(32'h684, 32'h0);
    mcoreClass.set_mregs(32'h685, 32'h0);
    mcoreClass.set_mregs(32'h686, 32'h0);
    mcoreClass.set_mregs(32'h687, 32'h0);
    mcoreClass.set_mregs(32'h688, 32'h0);
    mcoreClass.set_mregs(32'h689, 32'h0);
    mcoreClass.set_mregs(32'h68a, 32'h0);
    mcoreClass.set_mregs(32'h68b, 32'h0);
    mcoreClass.set_mregs(32'h68c, 32'h0);
    mcoreClass.set_mregs(32'h68d, 32'h0);
    mcoreClass.set_mregs(32'h68e, 32'h0);
    mcoreClass.set_mregs(32'h68f, 32'h0);
    mcoreClass.set_mregs(32'h690, 32'h0);
    mcoreClass.set_mregs(32'h691, 32'h0);
    mcoreClass.set_mregs(32'h692, 32'h0);
    mcoreClass.set_mregs(32'h693, 32'h0);
    mcoreClass.set_mregs(32'h694, 32'h0);
    mcoreClass.set_mregs(32'h695, 32'h0);
    mcoreClass.set_mregs(32'h696, 32'h0);
    mcoreClass.set_mregs(32'h697, 32'h0);
    mcoreClass.set_mregs(32'h698, 32'h0);
    mcoreClass.set_mregs(32'h699, 32'h0);
    mcoreClass.set_mregs(32'h69a, 32'h0);
    mcoreClass.set_mregs(32'h69b, 32'h0);
    mcoreClass.set_mregs(32'h69c, 32'h0);
    mcoreClass.set_mregs(32'h69d, 32'h0);
    mcoreClass.set_mregs(32'h69e, 32'h0);
    mcoreClass.set_mregs(32'h69f, 32'h0);
    mcoreClass.set_mregs(32'h6a0, 32'h0);
    mcoreClass.set_mregs(32'h6a1, 32'h0);
    mcoreClass.set_mregs(32'h6a2, 32'h0);
    mcoreClass.set_mregs(32'h6a3, 32'h0);
    mcoreClass.set_mregs(32'h6a4, 32'h0);
    mcoreClass.set_mregs(32'h6a5, 32'h0);
    mcoreClass.set_mregs(32'h6a6, 32'h0);
    mcoreClass.set_mregs(32'h6a7, 32'h0);
    mcoreClass.set_mregs(32'h6a8, 32'h0);
    mcoreClass.set_mregs(32'h6a9, 32'h0);
    mcoreClass.set_mregs(32'h6aa, 32'h0);
    mcoreClass.set_mregs(32'h6ab, 32'h0);
    mcoreClass.set_mregs(32'h6ac, 32'h0);
    mcoreClass.set_mregs(32'h6ad, 32'h0);
    mcoreClass.set_mregs(32'h6ae, 32'h0);
    mcoreClass.set_mregs(32'h6af, 32'h0);
    mcoreClass.set_mregs(32'h6b0, 32'h0);
    mcoreClass.set_mregs(32'h6b1, 32'h0);
    mcoreClass.set_mregs(32'h6b2, 32'h0);
    mcoreClass.set_mregs(32'h6b3, 32'h0);
    mcoreClass.set_mregs(32'h6b4, 32'h0);
    mcoreClass.set_mregs(32'h6b5, 32'h0);
    mcoreClass.set_mregs(32'h6b6, 32'h0);
    mcoreClass.set_mregs(32'h6b7, 32'h0);
    mcoreClass.set_mregs(32'h6b8, 32'h0);
    mcoreClass.set_mregs(32'h6b9, 32'h0);
    mcoreClass.set_mregs(32'h6ba, 32'h0);
    mcoreClass.set_mregs(32'h6bb, 32'h0);
    mcoreClass.set_mregs(32'h6bc, 32'h0);
    mcoreClass.set_mregs(32'h6bd, 32'h0);
    mcoreClass.set_mregs(32'h6be, 32'h0);
    mcoreClass.set_mregs(32'h6bf, 32'h0);
    mcoreClass.set_mregs(32'h6c0, 32'h0);
    mcoreClass.set_mregs(32'h6c1, 32'h0);
    mcoreClass.set_mregs(32'h6c2, 32'h0);
    mcoreClass.set_mregs(32'h6c3, 32'h0);
    mcoreClass.set_mregs(32'h6c4, 32'h0);
    mcoreClass.set_mregs(32'h6c5, 32'h0);
    mcoreClass.set_mregs(32'h6c6, 32'h0);
    mcoreClass.set_mregs(32'h6c7, 32'h0);
    mcoreClass.set_mregs(32'h6c8, 32'h0);
    mcoreClass.set_mregs(32'h6c9, 32'h0);
    mcoreClass.set_mregs(32'h6ca, 32'h0);
    mcoreClass.set_mregs(32'h6cb, 32'h0);
    mcoreClass.set_mregs(32'h6cc, 32'h0);
    mcoreClass.set_mregs(32'h6cd, 32'h0);
    mcoreClass.set_mregs(32'h6ce, 32'h0);
    mcoreClass.set_mregs(32'h6cf, 32'h0);
    mcoreClass.set_mregs(32'h6d0, 32'h0);
    mcoreClass.set_mregs(32'h6d1, 32'h0);
    mcoreClass.set_mregs(32'h6d2, 32'h0);
    mcoreClass.set_mregs(32'h6d3, 32'h0);
    mcoreClass.set_mregs(32'h6d4, 32'h0);
    mcoreClass.set_mregs(32'h6d5, 32'h0);
    mcoreClass.set_mregs(32'h6d6, 32'h0);
    mcoreClass.set_mregs(32'h6d7, 32'h0);
    mcoreClass.set_mregs(32'h6d8, 32'h0);
    mcoreClass.set_mregs(32'h6d9, 32'h0);
    mcoreClass.set_mregs(32'h6da, 32'h0);
    mcoreClass.set_mregs(32'h6db, 32'h0);
    mcoreClass.set_mregs(32'h6dc, 32'h0);
    mcoreClass.set_mregs(32'h6dd, 32'h0);
    mcoreClass.set_mregs(32'h6de, 32'h0);
    mcoreClass.set_mregs(32'h6df, 32'h0);
    mcoreClass.set_mregs(32'h6e0, 32'h0);
    mcoreClass.set_mregs(32'h6e1, 32'h0);
    mcoreClass.set_mregs(32'h6e2, 32'h0);
    mcoreClass.set_mregs(32'h6e3, 32'h0);
    mcoreClass.set_mregs(32'h6e4, 32'h0);
    mcoreClass.set_mregs(32'h6e5, 32'h0);
    mcoreClass.set_mregs(32'h6e6, 32'h0);
    mcoreClass.set_mregs(32'h6e7, 32'h0);
    mcoreClass.set_mregs(32'h6e8, 32'h0);
    mcoreClass.set_mregs(32'h6e9, 32'h0);
    mcoreClass.set_mregs(32'h6ea, 32'h0);
    mcoreClass.set_mregs(32'h6eb, 32'h0);
    mcoreClass.set_mregs(32'h6ec, 32'h0);
    mcoreClass.set_mregs(32'h6ed, 32'h0);
    mcoreClass.set_mregs(32'h6ee, 32'h0);
    mcoreClass.set_mregs(32'h6ef, 32'h0);
    mcoreClass.set_mregs(32'h6f0, 32'h0);
    mcoreClass.set_mregs(32'h6f1, 32'h0);
    mcoreClass.set_mregs(32'h6f2, 32'h0);
    mcoreClass.set_mregs(32'h6f3, 32'h0);
    mcoreClass.set_mregs(32'h6f4, 32'h0);
    mcoreClass.set_mregs(32'h6f5, 32'h0);
    mcoreClass.set_mregs(32'h6f6, 32'h0);
    mcoreClass.set_mregs(32'h6f7, 32'h0);
    mcoreClass.set_mregs(32'h6f8, 32'h0);
    mcoreClass.set_mregs(32'h6f9, 32'h0);
    mcoreClass.set_mregs(32'h6fa, 32'h0);
    mcoreClass.set_mregs(32'h6fb, 32'h0);
    mcoreClass.set_mregs(32'h6fc, 32'h0);
    mcoreClass.set_mregs(32'h6fd, 32'h0);
    mcoreClass.set_mregs(32'h6fe, 32'h0);
    mcoreClass.set_mregs(32'h6ff, 32'h0);
    mcoreClass.set_mregs(32'h700, 32'h0);
    mcoreClass.set_mregs(32'h701, 32'h0);
    mcoreClass.set_mregs(32'h702, 32'h0);
    mcoreClass.set_mregs(32'h703, 32'h0);
    mcoreClass.set_mregs(32'h704, 32'h0);
    mcoreClass.set_mregs(32'h705, 32'h0);
    mcoreClass.set_mregs(32'h706, 32'h0);
    mcoreClass.set_mregs(32'h707, 32'h0);
    mcoreClass.set_mregs(32'h708, 32'h0);
    mcoreClass.set_mregs(32'h709, 32'h0);
    mcoreClass.set_mregs(32'h70a, 32'h0);
    mcoreClass.set_mregs(32'h70b, 32'h0);
    mcoreClass.set_mregs(32'h70c, 32'h0);
    mcoreClass.set_mregs(32'h70d, 32'h0);
    mcoreClass.set_mregs(32'h70e, 32'h0);
    mcoreClass.set_mregs(32'h70f, 32'h0);
    mcoreClass.set_mregs(32'h710, 32'h0);
    mcoreClass.set_mregs(32'h711, 32'h0);
    mcoreClass.set_mregs(32'h712, 32'h0);
    mcoreClass.set_mregs(32'h713, 32'h0);
    mcoreClass.set_mregs(32'h714, 32'h0);
    mcoreClass.set_mregs(32'h715, 32'h0);
    mcoreClass.set_mregs(32'h716, 32'h0);
    mcoreClass.set_mregs(32'h717, 32'h0);
    mcoreClass.set_mregs(32'h718, 32'h0);
    mcoreClass.set_mregs(32'h719, 32'h0);
    mcoreClass.set_mregs(32'h71a, 32'h0);
    mcoreClass.set_mregs(32'h71b, 32'h0);
    mcoreClass.set_mregs(32'h71c, 32'h0);
    mcoreClass.set_mregs(32'h71d, 32'h0);
    mcoreClass.set_mregs(32'h71e, 32'h0);
    mcoreClass.set_mregs(32'h71f, 32'h0);
    mcoreClass.set_mregs(32'h720, 32'h0);
    mcoreClass.set_mregs(32'h721, 32'h0);
    mcoreClass.set_mregs(32'h722, 32'h0);
    mcoreClass.set_mregs(32'h723, 32'h0);
    mcoreClass.set_mregs(32'h724, 32'h0);
    mcoreClass.set_mregs(32'h725, 32'h0);
    mcoreClass.set_mregs(32'h726, 32'h0);
    mcoreClass.set_mregs(32'h727, 32'h0);
    mcoreClass.set_mregs(32'h728, 32'h0);
    mcoreClass.set_mregs(32'h729, 32'h0);
    mcoreClass.set_mregs(32'h72a, 32'h0);
    mcoreClass.set_mregs(32'h72b, 32'h0);
    mcoreClass.set_mregs(32'h72c, 32'h0);
    mcoreClass.set_mregs(32'h72d, 32'h0);
    mcoreClass.set_mregs(32'h72e, 32'h0);
    mcoreClass.set_mregs(32'h72f, 32'h0);
    mcoreClass.set_mregs(32'h730, 32'h0);
    mcoreClass.set_mregs(32'h731, 32'h0);
    mcoreClass.set_mregs(32'h732, 32'h0);
    mcoreClass.set_mregs(32'h733, 32'h0);
    mcoreClass.set_mregs(32'h734, 32'h0);
    mcoreClass.set_mregs(32'h735, 32'h0);
    mcoreClass.set_mregs(32'h736, 32'h0);
    mcoreClass.set_mregs(32'h737, 32'h0);
    mcoreClass.set_mregs(32'h738, 32'h0);
    mcoreClass.set_mregs(32'h739, 32'h0);
    mcoreClass.set_mregs(32'h73a, 32'h0);
    mcoreClass.set_mregs(32'h73b, 32'h0);
    mcoreClass.set_mregs(32'h73c, 32'h0);
    mcoreClass.set_mregs(32'h73d, 32'h0);
    mcoreClass.set_mregs(32'h73e, 32'h0);
    mcoreClass.set_mregs(32'h73f, 32'h0);
    mcoreClass.set_mregs(32'h740, 32'h0);
    mcoreClass.set_mregs(32'h741, 32'h0);
    mcoreClass.set_mregs(32'h742, 32'h0);
    mcoreClass.set_mregs(32'h743, 32'h0);
    mcoreClass.set_mregs(32'h744, 32'h0);
    mcoreClass.set_mregs(32'h745, 32'h0);
    mcoreClass.set_mregs(32'h746, 32'h0);
    mcoreClass.set_mregs(32'h747, 32'h0);
    mcoreClass.set_mregs(32'h748, 32'h0);
    mcoreClass.set_mregs(32'h749, 32'h0);
    mcoreClass.set_mregs(32'h74a, 32'h0);
    mcoreClass.set_mregs(32'h74b, 32'h0);
    mcoreClass.set_mregs(32'h74c, 32'h0);
    mcoreClass.set_mregs(32'h74d, 32'h0);
    mcoreClass.set_mregs(32'h74e, 32'h0);
    mcoreClass.set_mregs(32'h74f, 32'h0);
    mcoreClass.set_mregs(32'h750, 32'h0);
    mcoreClass.set_mregs(32'h751, 32'h0);
    mcoreClass.set_mregs(32'h752, 32'h0);
    mcoreClass.set_mregs(32'h753, 32'h0);
    mcoreClass.set_mregs(32'h754, 32'h0);
    mcoreClass.set_mregs(32'h755, 32'h0);
    mcoreClass.set_mregs(32'h756, 32'h0);
    mcoreClass.set_mregs(32'h757, 32'h0);
    mcoreClass.set_mregs(32'h758, 32'h0);
    mcoreClass.set_mregs(32'h759, 32'h0);
    mcoreClass.set_mregs(32'h75a, 32'h0);
    mcoreClass.set_mregs(32'h75b, 32'h0);
    mcoreClass.set_mregs(32'h75c, 32'h0);
    mcoreClass.set_mregs(32'h75d, 32'h0);
    mcoreClass.set_mregs(32'h75e, 32'h0);
    mcoreClass.set_mregs(32'h75f, 32'h0);
    mcoreClass.set_mregs(32'h760, 32'h0);
    mcoreClass.set_mregs(32'h761, 32'h0);
    mcoreClass.set_mregs(32'h762, 32'h0);
    mcoreClass.set_mregs(32'h763, 32'h0);
    mcoreClass.set_mregs(32'h764, 32'h0);
    mcoreClass.set_mregs(32'h765, 32'h0);
    mcoreClass.set_mregs(32'h766, 32'h0);
    mcoreClass.set_mregs(32'h767, 32'h0);
    mcoreClass.set_mregs(32'h768, 32'h0);
    mcoreClass.set_mregs(32'h769, 32'h0);
    mcoreClass.set_mregs(32'h76a, 32'h0);
    mcoreClass.set_mregs(32'h76b, 32'h0);
    mcoreClass.set_mregs(32'h76c, 32'h0);
    mcoreClass.set_mregs(32'h76d, 32'h0);
    mcoreClass.set_mregs(32'h76e, 32'h0);
    mcoreClass.set_mregs(32'h76f, 32'h0);
    mcoreClass.set_mregs(32'h770, 32'h0);
    mcoreClass.set_mregs(32'h771, 32'h0);
    mcoreClass.set_mregs(32'h772, 32'h0);
    mcoreClass.set_mregs(32'h773, 32'h0);
    mcoreClass.set_mregs(32'h774, 32'h0);
    mcoreClass.set_mregs(32'h775, 32'h0);
    mcoreClass.set_mregs(32'h776, 32'h0);
    mcoreClass.set_mregs(32'h777, 32'h0);
    mcoreClass.set_mregs(32'h778, 32'h0);
    mcoreClass.set_mregs(32'h779, 32'h0);
    mcoreClass.set_mregs(32'h77a, 32'h0);
    mcoreClass.set_mregs(32'h77b, 32'h0);
    mcoreClass.set_mregs(32'h77c, 32'h0);
    mcoreClass.set_mregs(32'h77d, 32'h0);
    mcoreClass.set_mregs(32'h77e, 32'h0);
    mcoreClass.set_mregs(32'h77f, 32'h0);
    mcoreClass.set_mregs(32'h780, 32'h0);
    mcoreClass.set_mregs(32'h781, 32'h0);
    mcoreClass.set_mregs(32'h782, 32'h0);
    mcoreClass.set_mregs(32'h783, 32'h0);
    mcoreClass.set_mregs(32'h784, 32'h0);
    mcoreClass.set_mregs(32'h785, 32'h0);
    mcoreClass.set_mregs(32'h786, 32'h0);
    mcoreClass.set_mregs(32'h787, 32'h0);
    mcoreClass.set_mregs(32'h788, 32'h0);
    mcoreClass.set_mregs(32'h789, 32'h0);
    mcoreClass.set_mregs(32'h78a, 32'h0);
    mcoreClass.set_mregs(32'h78b, 32'h0);
    mcoreClass.set_mregs(32'h78c, 32'h0);
    mcoreClass.set_mregs(32'h78d, 32'h0);
    mcoreClass.set_mregs(32'h78e, 32'h0);
    mcoreClass.set_mregs(32'h78f, 32'h0);
    mcoreClass.set_mregs(32'h790, 32'h0);
    mcoreClass.set_mregs(32'h791, 32'h0);
    mcoreClass.set_mregs(32'h792, 32'h0);
    mcoreClass.set_mregs(32'h793, 32'h0);
    mcoreClass.set_mregs(32'h794, 32'h0);
    mcoreClass.set_mregs(32'h795, 32'h0);
    mcoreClass.set_mregs(32'h796, 32'h0);
    mcoreClass.set_mregs(32'h797, 32'h0);
    mcoreClass.set_mregs(32'h798, 32'h0);
    mcoreClass.set_mregs(32'h799, 32'h0);
    mcoreClass.set_mregs(32'h79a, 32'h0);
    mcoreClass.set_mregs(32'h79b, 32'h0);
    mcoreClass.set_mregs(32'h79c, 32'h0);
    mcoreClass.set_mregs(32'h79d, 32'h0);
    mcoreClass.set_mregs(32'h79e, 32'h0);
    mcoreClass.set_mregs(32'h79f, 32'h0);
    mcoreClass.set_mregs(32'h7a0, 32'h0);
    mcoreClass.set_mregs(32'h7a1, 32'h0);
    mcoreClass.set_mregs(32'h7a2, 32'h0);
    mcoreClass.set_mregs(32'h7a3, 32'h0);
    mcoreClass.set_mregs(32'h7a4, 32'h0);
    mcoreClass.set_mregs(32'h7a5, 32'h0);
    mcoreClass.set_mregs(32'h7a6, 32'h0);
    mcoreClass.set_mregs(32'h7a7, 32'h0);
    mcoreClass.set_mregs(32'h7a8, 32'h0);
    mcoreClass.set_mregs(32'h7a9, 32'h0);
    mcoreClass.set_mregs(32'h7aa, 32'h0);
    mcoreClass.set_mregs(32'h7ab, 32'h0);
    mcoreClass.set_mregs(32'h7ac, 32'h0);
    mcoreClass.set_mregs(32'h7ad, 32'h0);
    mcoreClass.set_mregs(32'h7ae, 32'h0);
    mcoreClass.set_mregs(32'h7af, 32'h0);
    mcoreClass.set_mregs(32'h7b0, 32'h0);
    mcoreClass.set_mregs(32'h7b1, 32'h0);
    mcoreClass.set_mregs(32'h7b2, 32'h0);
    mcoreClass.set_mregs(32'h7b3, 32'h0);
    mcoreClass.set_mregs(32'h7b4, 32'h0);
    mcoreClass.set_mregs(32'h7b5, 32'h0);
    mcoreClass.set_mregs(32'h7b6, 32'h0);
    mcoreClass.set_mregs(32'h7b7, 32'h0);
    mcoreClass.set_mregs(32'h7b8, 32'h0);
    mcoreClass.set_mregs(32'h7b9, 32'h0);
    mcoreClass.set_mregs(32'h7ba, 32'h0);
    mcoreClass.set_mregs(32'h7bb, 32'h0);
    mcoreClass.set_mregs(32'h7bc, 32'h0);
    mcoreClass.set_mregs(32'h7bd, 32'h0);
    mcoreClass.set_mregs(32'h7be, 32'h0);
    mcoreClass.set_mregs(32'h7bf, 32'h0);
    mcoreClass.set_mregs(32'h7c0, 32'h0);
    mcoreClass.set_mregs(32'h7c1, 32'h0);
    mcoreClass.set_mregs(32'h7c2, 32'h0);
    mcoreClass.set_mregs(32'h7c3, 32'h0);
    mcoreClass.set_mregs(32'h7c4, 32'h0);
    mcoreClass.set_mregs(32'h7c5, 32'h0);
    mcoreClass.set_mregs(32'h7c6, 32'h0);
    mcoreClass.set_mregs(32'h7c7, 32'h0);
    mcoreClass.set_mregs(32'h7c8, 32'h0);
    mcoreClass.set_mregs(32'h7c9, 32'h0);
    mcoreClass.set_mregs(32'h7ca, 32'h0);
    mcoreClass.set_mregs(32'h7cb, 32'h0);
    mcoreClass.set_mregs(32'h7cc, 32'h0);
    mcoreClass.set_mregs(32'h7cd, 32'h0);
    mcoreClass.set_mregs(32'h7ce, 32'h0);
    mcoreClass.set_mregs(32'h7cf, 32'h0);
    mcoreClass.set_mregs(32'h7d0, 32'h0);
    mcoreClass.set_mregs(32'h7d1, 32'h0);
    mcoreClass.set_mregs(32'h7d2, 32'h0);
    mcoreClass.set_mregs(32'h7d3, 32'h0);
    mcoreClass.set_mregs(32'h7d4, 32'h0);
    mcoreClass.set_mregs(32'h7d5, 32'h0);
    mcoreClass.set_mregs(32'h7d6, 32'h0);
    mcoreClass.set_mregs(32'h7d7, 32'h0);
    mcoreClass.set_mregs(32'h7d8, 32'h0);
    mcoreClass.set_mregs(32'h7d9, 32'h0);
    mcoreClass.set_mregs(32'h7da, 32'h0);
    mcoreClass.set_mregs(32'h7db, 32'h0);
    mcoreClass.set_mregs(32'h7dc, 32'h0);
    mcoreClass.set_mregs(32'h7dd, 32'h0);
    mcoreClass.set_mregs(32'h7de, 32'h0);
    mcoreClass.set_mregs(32'h7df, 32'h0);
    mcoreClass.set_mregs(32'h7e0, 32'h0);
    mcoreClass.set_mregs(32'h7e1, 32'h0);
    mcoreClass.set_mregs(32'h7e2, 32'h0);
    mcoreClass.set_mregs(32'h7e3, 32'h0);
    mcoreClass.set_mregs(32'h7e4, 32'h0);
    mcoreClass.set_mregs(32'h7e5, 32'h0);
    mcoreClass.set_mregs(32'h7e6, 32'h0);
    mcoreClass.set_mregs(32'h7e7, 32'h0);
    mcoreClass.set_mregs(32'h7e8, 32'h0);
    mcoreClass.set_mregs(32'h7e9, 32'h0);
    mcoreClass.set_mregs(32'h7ea, 32'h0);
    mcoreClass.set_mregs(32'h7eb, 32'h0);
    mcoreClass.set_mregs(32'h7ec, 32'h0);
    mcoreClass.set_mregs(32'h7ed, 32'h0);
    mcoreClass.set_mregs(32'h7ee, 32'h0);
    mcoreClass.set_mregs(32'h7ef, 32'h0);
    mcoreClass.set_mregs(32'h7f0, 32'h65);
    mcoreClass.set_mregs(32'h7f1, 32'h0);
    mcoreClass.set_mregs(32'h7f2, 32'h0);
    mcoreClass.set_mregs(32'h7f3, 32'h0);
    mcoreClass.set_mregs(32'h7f4, 32'hffffffff);
    mcoreClass.set_mregs(32'h7f5, 32'h0);
    mcoreClass.set_mregs(32'h7f6, 32'h0);
    mcoreClass.set_mregs(32'h7f7, 32'h0);
    mcoreClass.set_mregs(32'h7f8, 32'h0);
    mcoreClass.set_mregs(32'h7f9, 32'h0);
    mcoreClass.set_mregs(32'h7fa, 32'h0);
    mcoreClass.set_mregs(32'h7fb, 32'h0);
    mcoreClass.set_mregs(32'h7fc, 32'h0);
    mcoreClass.set_mregs(32'h7fd, 32'h0);
    mcoreClass.set_mregs(32'h7fe, 32'h0);
    mcoreClass.set_mregs(32'h7ff, 32'h0);
    mcoreClass.set_wmod(32'h500);


/*Setup mregs end*/
/*Setup PDEC begin*/
    mcoreClass.set_utils_reg(32'h20, 32'h0);
    mcoreClass.set_utils_reg(32'h21, 32'hf);
    mcoreClass.set_utils_reg(32'h22, 32'h1);
/*Setup PDEC end*/
    mcoreClass.load_plut(PLUT);
endtask

